`timescale 1ns/1ps
`default_nettype none

module fpga_agc(p4VDC, p4VSW, GND, SIM_RST, SIM_CLK, BLKUPL_n, BMGXM, BMGXP, BMGYM, BMGYP, BMGZM, BMGZP, CAURST, CDUFAL, CDUXM, CDUXP, CDUYM, CDUYP, CDUZM, CDUZP, CLOCK, CTLSAT, DBLTST, DKBSNC, DKEND, DKSTRT, DOSCAL, FLTOUT, FREFUN, GATEX_n, GATEY_n, GATEZ_n, GCAPCL, GUIREL, HOLFUN, IMUCAG, IMUFAL, IMUOPR, IN3008, IN3212, IN3213, IN3214, IN3216, IN3301, ISSTOR, LEMATT, LFTOFF, LRIN0, LRIN1, LRRLSC, LVDAGD, MAINRS, MAMU, MANmP, MANmR, MANmY, MANpP, MANpR, MANpY, MARK, MDT01, MDT02, MDT03, MDT04, MDT05, MDT06, MDT07, MDT08, MDT09, MDT10, MDT11, MDT12, MDT13, MDT14, MDT15, MDT16, MKEY1, MKEY2, MKEY3, MKEY4, MKEY5, MLDCH, MLOAD, MNHNC, MNHRPT, MNHSBF, MNIMmP, MNIMmR, MNIMmY, MNIMpP, MNIMpR, MNIMpY, MONPAR, MONWBK, MRDCH, MREAD, MRKREJ, MRKRST, MSTP, MSTRT, MTCSAI, MYCLMP, NAVRST, NHALGA, NHVFAL, NKEY1, NKEY2, NKEY3, NKEY4, NKEY5, OPCDFL, OPMSW2, OPMSW3, PCHGOF, PIPAXm, PIPAXp, PIPAYm, PIPAYp, PIPAZm, PIPAZp, ROLGOF, RRIN0, RRIN1, RRPONA, RRRLSC, S4BSAB, SBYBUT, SCAFAL, SHAFTM, SHAFTP, SIGNX, SIGNY, SIGNZ, SMSEPR, SPSRDY, STRPRS, STRT2, TEMPIN, TRANmX, TRANmY, TRANmZ, TRANpX, TRANpY, TRANpZ, TRNM, TRNP, TRST10, TRST9, ULLTHR, UPL0, UPL1, VFAIL, XLNK0, XLNK1, ZEROP, n2FSFAL, CDUXDM, CDUXDP, CDUYDM, CDUYDP, CDUZDM, CDUZDP, CLK, COMACT, DKDATA, ELSNCM, ELSNCN, KYRLS, MBR1, MBR2, MCTRAL_n, MGOJAM, MGP_n, MIIP, MINHL, MINKL, MNISQ, MON800, MONWT, MOSCAL_n, MPAL_n, MPIPAL_n, MRAG, MRCH, MREQIN, MRGG, MRLG, MRPTAL_n, MRSC, MRULOG, MSCAFL_n, MSCDBL_n, MSP, MSQ10, MSQ11, MSQ12, MSQ13, MSQ14, MSQ16, MSQEXT, MST1, MST2, MST3, MSTPIT_n, MT01, MT02, MT03, MT04, MT05, MT06, MT07, MT08, MT09, MT10, MT11, MT12, MTCAL_n, MTCSA_n, MVFAIL_n, MWAG, MWARNF_n, MWATCH_n, MWBBEG, MWBG, MWCH, MWEBG, MWFBG, MWG, MWL01, MWL02, MWL03, MWL04, MWL05, MWL06, MWL07, MWL08, MWL09, MWL10, MWL11, MWL12, MWL13, MWL14, MWL15, MWL16, MWLG, MWQG, MWSG, MWYG, MWZG, OPEROR, OUTCOM, PIPASW, PIPDAT, RESTRT, RLYB01, RLYB02, RLYB03, RLYB04, RLYB05, RLYB06, RLYB07, RLYB08, RLYB09, RLYB10, RLYB11, RYWD12, RYWD13, RYWD14, RYWD16, SBYLIT, SBYREL_n, TMPCAU, UPLACT, VNFLSH);
    input wire p4VDC;
    input wire p4VSW;
    input wire GND;
    input wire SIM_RST;
    input wire SIM_CLK;
    input wire BLKUPL_n;
    input wire BMGXM;
    input wire BMGXP;
    input wire BMGYM;
    input wire BMGYP;
    input wire BMGZM;
    input wire BMGZP;
    input wire CAURST;
    input wire CDUFAL;
    input wire CDUXM;
    input wire CDUXP;
    input wire CDUYM;
    input wire CDUYP;
    input wire CDUZM;
    input wire CDUZP;
    input wire CLOCK;
    input wire CTLSAT;
    input wire DBLTST;
    input wire DKBSNC;
    input wire DKEND;
    input wire DKSTRT;
    input wire DOSCAL;
    input wire FLTOUT;
    input wire FREFUN;
    input wire GATEX_n;
    input wire GATEY_n;
    input wire GATEZ_n;
    input wire GCAPCL;
    input wire GUIREL;
    input wire HOLFUN;
    input wire IMUCAG;
    input wire IMUFAL;
    input wire IMUOPR;
    input wire IN3008;
    input wire IN3212;
    input wire IN3213;
    input wire IN3214;
    input wire IN3216;
    input wire IN3301;
    input wire ISSTOR;
    input wire LEMATT;
    input wire LFTOFF;
    input wire LRIN0;
    input wire LRIN1;
    input wire LRRLSC;
    input wire LVDAGD;
    input wire MAINRS;
    input wire MAMU;
    input wire MANmP;
    input wire MANmR;
    input wire MANmY;
    input wire MANpP;
    input wire MANpR;
    input wire MANpY;
    input wire MARK;
    input wire MDT01;
    input wire MDT02;
    input wire MDT03;
    input wire MDT04;
    input wire MDT05;
    input wire MDT06;
    input wire MDT07;
    input wire MDT08;
    input wire MDT09;
    input wire MDT10;
    input wire MDT11;
    input wire MDT12;
    input wire MDT13;
    input wire MDT14;
    input wire MDT15;
    input wire MDT16;
    input wire MKEY1;
    input wire MKEY2;
    input wire MKEY3;
    input wire MKEY4;
    input wire MKEY5;
    input wire MLDCH;
    input wire MLOAD;
    input wire MNHNC;
    input wire MNHRPT;
    input wire MNHSBF;
    input wire MNIMmP;
    input wire MNIMmR;
    input wire MNIMmY;
    input wire MNIMpP;
    input wire MNIMpR;
    input wire MNIMpY;
    input wire MONPAR;
    input wire MONWBK;
    input wire MRDCH;
    input wire MREAD;
    input wire MRKREJ;
    input wire MRKRST;
    input wire MSTP;
    input wire MSTRT;
    input wire MTCSAI;
    input wire MYCLMP;
    input wire NAVRST;
    input wire NHALGA;
    input wire NHVFAL;
    input wire NKEY1;
    input wire NKEY2;
    input wire NKEY3;
    input wire NKEY4;
    input wire NKEY5;
    input wire OPCDFL;
    input wire OPMSW2;
    input wire OPMSW3;
    input wire PCHGOF;
    input wire PIPAXm;
    input wire PIPAXp;
    input wire PIPAYm;
    input wire PIPAYp;
    input wire PIPAZm;
    input wire PIPAZp;
    input wire ROLGOF;
    input wire RRIN0;
    input wire RRIN1;
    input wire RRPONA;
    input wire RRRLSC;
    input wire S4BSAB;
    input wire SBYBUT;
    input wire SCAFAL;
    input wire SHAFTM;
    input wire SHAFTP;
    input wire SIGNX;
    input wire SIGNY;
    input wire SIGNZ;
    input wire SMSEPR;
    input wire SPSRDY;
    input wire STRPRS;
    input wire STRT2;
    input wire TEMPIN;
    input wire TRANmX;
    input wire TRANmY;
    input wire TRANmZ;
    input wire TRANpX;
    input wire TRANpY;
    input wire TRANpZ;
    input wire TRNM;
    input wire TRNP;
    input wire TRST10;
    input wire TRST9;
    input wire ULLTHR;
    input wire UPL0;
    input wire UPL1;
    input wire VFAIL;
    input wire XLNK0;
    input wire XLNK1;
    input wire ZEROP;
    input wire n2FSFAL;
    output wire CDUXDM;
    output wire CDUXDP;
    output wire CDUYDM;
    output wire CDUYDP;
    output wire CDUZDM;
    output wire CDUZDP;
    output wire CLK;
    output wire COMACT;
    output wire DKDATA;
    output wire ELSNCM;
    output wire ELSNCN;
    output wire KYRLS;
    output wire MBR1;
    output wire MBR2;
    output wire MCTRAL_n;
    output wire MGOJAM;
    output wire MGP_n;
    output wire MIIP;
    output wire MINHL;
    output wire MINKL;
    output wire MNISQ;
    output wire MON800;
    output wire MONWT;
    output wire MOSCAL_n;
    output wire MPAL_n;
    output wire MPIPAL_n;
    output wire MRAG;
    output wire MRCH;
    output wire MREQIN;
    output wire MRGG;
    output wire MRLG;
    output wire MRPTAL_n;
    output wire MRSC;
    output wire MRULOG;
    output wire MSCAFL_n;
    output wire MSCDBL_n;
    output wire MSP;
    output wire MSQ10;
    output wire MSQ11;
    output wire MSQ12;
    output wire MSQ13;
    output wire MSQ14;
    output wire MSQ16;
    output wire MSQEXT;
    output wire MST1;
    output wire MST2;
    output wire MST3;
    output wire MSTPIT_n;
    output wire MT01;
    output wire MT02;
    output wire MT03;
    output wire MT04;
    output wire MT05;
    output wire MT06;
    output wire MT07;
    output wire MT08;
    output wire MT09;
    output wire MT10;
    output wire MT11;
    output wire MT12;
    output wire MTCAL_n;
    output wire MTCSA_n;
    output wire MVFAIL_n;
    output wire MWAG;
    output wire MWARNF_n;
    output wire MWATCH_n;
    output wire MWBBEG;
    output wire MWBG;
    output wire MWCH;
    output wire MWEBG;
    output wire MWFBG;
    output wire MWG;
    output wire MWL01;
    output wire MWL02;
    output wire MWL03;
    output wire MWL04;
    output wire MWL05;
    output wire MWL06;
    output wire MWL07;
    output wire MWL08;
    output wire MWL09;
    output wire MWL10;
    output wire MWL11;
    output wire MWL12;
    output wire MWL13;
    output wire MWL14;
    output wire MWL15;
    output wire MWL16;
    output wire MWLG;
    output wire MWQG;
    output wire MWSG;
    output wire MWYG;
    output wire MWZG;
    output wire OPEROR;
    output wire OUTCOM;
    output wire PIPASW;
    output wire PIPDAT;
    output wire RESTRT;
    output wire RLYB01;
    output wire RLYB02;
    output wire RLYB03;
    output wire RLYB04;
    output wire RLYB05;
    output wire RLYB06;
    output wire RLYB07;
    output wire RLYB08;
    output wire RLYB09;
    output wire RLYB10;
    output wire RLYB11;
    output wire RYWD12;
    output wire RYWD13;
    output wire RYWD14;
    output wire RYWD16;
    output wire SBYLIT;
    output wire SBYREL_n;
    output wire TMPCAU;
    output wire UPLACT;
    output wire VNFLSH;
    wire A15_n;
    wire A16_n;
    wire A2XG_n;
    wire A2X_n;
    wire A2X_n_U5012_10;
    wire A2X_n_U5044_8;
    wire A2X_n_U6004_6;
    wire AD0;
    wire ADS0;
    wire AGCWAR;
    wire ALGA;
    wire ALTEST;
    wire ALTM;
    wire AUG0_n;
    wire B15X;
    wire BKTF_n;
    wire BMAGXM;
    wire BMAGXP;
    wire BMAGYM;
    wire BMAGYP;
    wire BMAGZM;
    wire BMAGZP;
    wire BR1;
    wire BR12B_n;
    wire BR1B2B;
    wire BR1B2B_n;
    wire BR1B2_n;
    wire BR1_n;
    wire BR2;
    wire BR2_n;
    wire BRDIF_n;
    wire BXVX;
    wire C24A;
    wire C25A;
    wire C26A;
    wire C27A;
    wire C30A;
    wire C31A;
    wire C32A;
    wire C32M;
    wire C32P;
    wire C33A;
    wire C33M;
    wire C33P;
    wire C34A;
    wire C34M;
    wire C34P;
    wire C35A;
    wire C35M;
    wire C35P;
    wire C36A;
    wire C36M;
    wire C36P;
    wire C37A;
    wire C37M;
    wire C37P;
    wire C40A;
    wire C40M;
    wire C40P;
    wire C41A;
    wire C41M;
    wire C41P;
    wire C45R;
    wire C50A;
    wire C51A;
    wire C52A;
    wire C53A;
    wire C54A;
    wire C55A;
    wire CA2_n;
    wire CA3_n;
    wire CA4_n;
    wire CA5_n;
    wire CA6_n;
    wire CAD1;
    wire CAD2;
    wire CAD3;
    wire CAD4;
    wire CAD5;
    wire CAD6;
    wire CAG;
    wire CBG;
    wire CCH11;
    wire CCH12;
    wire CCH13;
    wire CCH14;
    wire CCH33;
    wire CCH34;
    wire CCH35;
    wire CCHG_n;
    wire CCS0;
    wire CCS0_n;
    wire CDUSTB_n;
    wire CDUXD;
    wire CDUYD;
    wire CDUZD;
    wire CEBG;
    wire CFBG;
    wire CG13;
    wire CG23;
    wire CG26;
    wire CGG;
    wire CGMC;
    wire CH01;
    wire CH02;
    wire CH03;
    wire CH04;
    wire CH05;
    wire CH06;
    wire CH07;
    wire CH0705;
    wire CH0706;
    wire CH0707;
    wire CH08;
    wire CH09;
    wire CH10;
    wire CH11;
    wire CH1108;
    wire CH1109;
    wire CH1110;
    wire CH1111;
    wire CH1112;
    wire CH1113;
    wire CH1114;
    wire CH1116;
    wire CH12;
    wire CH1208;
    wire CH1209;
    wire CH1210;
    wire CH1211;
    wire CH1212;
    wire CH1213;
    wire CH1214;
    wire CH1216;
    wire CH13;
    wire CH1301;
    wire CH1302;
    wire CH1303;
    wire CH1304;
    wire CH1305;
    wire CH1306;
    wire CH1307;
    wire CH1308;
    wire CH1309;
    wire CH1310;
    wire CH1311;
    wire CH1316;
    wire CH14;
    wire CH1401;
    wire CH1402;
    wire CH1403;
    wire CH1404;
    wire CH1405;
    wire CH1406;
    wire CH1407;
    wire CH1408;
    wire CH1409;
    wire CH1410;
    wire CH1411;
    wire CH1412;
    wire CH1413;
    wire CH1414;
    wire CH1416;
    wire CH1501;
    wire CH1502;
    wire CH1503;
    wire CH1504;
    wire CH1505;
    wire CH16;
    wire CH1601;
    wire CH1602;
    wire CH1603;
    wire CH1604;
    wire CH1605;
    wire CH1606;
    wire CH1607;
    wire CH3201;
    wire CH3202;
    wire CH3203;
    wire CH3204;
    wire CH3205;
    wire CH3206;
    wire CH3207;
    wire CH3208;
    wire CH3209;
    wire CH3210;
    wire CH3310;
    wire CH3311;
    wire CH3312;
    wire CH3313;
    wire CH3314;
    wire CH3316;
    wire CHAT01;
    wire CHAT02;
    wire CHAT03;
    wire CHAT04;
    wire CHAT05;
    wire CHAT06;
    wire CHAT07;
    wire CHAT08;
    wire CHAT09;
    wire CHAT10;
    wire CHAT11;
    wire CHAT12;
    wire CHAT13;
    wire CHAT14;
    wire CHBT01;
    wire CHBT02;
    wire CHBT03;
    wire CHBT04;
    wire CHBT05;
    wire CHBT06;
    wire CHBT07;
    wire CHBT08;
    wire CHBT09;
    wire CHBT10;
    wire CHBT11;
    wire CHBT12;
    wire CHBT13;
    wire CHBT14;
    wire CHINC;
    wire CHINC_n;
    wire CHOR01_n;
    wire CHOR01_n_U16004_2;
    wire CHOR01_n_U16021_6;
    wire CHOR01_n_U17003_2;
    wire CHOR01_n_U17027_10;
    wire CHOR01_n_U24011_2;
    wire CHOR02_n;
    wire CHOR02_n_U16004_4;
    wire CHOR02_n_U16021_8;
    wire CHOR02_n_U17003_4;
    wire CHOR02_n_U17041_2;
    wire CHOR02_n_U24011_4;
    wire CHOR03_n;
    wire CHOR03_n_U16004_6;
    wire CHOR03_n_U16021_10;
    wire CHOR03_n_U17003_6;
    wire CHOR03_n_U17041_4;
    wire CHOR03_n_U24011_6;
    wire CHOR04_n;
    wire CHOR04_n_U16004_8;
    wire CHOR04_n_U16021_12;
    wire CHOR04_n_U17003_8;
    wire CHOR04_n_U17041_6;
    wire CHOR04_n_U24011_8;
    wire CHOR05_n;
    wire CHOR05_n_U16004_10;
    wire CHOR05_n_U16044_2;
    wire CHOR05_n_U17003_10;
    wire CHOR05_n_U17041_8;
    wire CHOR05_n_U24011_10;
    wire CHOR06_n;
    wire CHOR06_n_U16004_12;
    wire CHOR06_n_U16044_4;
    wire CHOR06_n_U17003_12;
    wire CHOR06_n_U17041_10;
    wire CHOR06_n_U24011_12;
    wire CHOR07_n;
    wire CHOR07_n_U16021_2;
    wire CHOR07_n_U16044_6;
    wire CHOR07_n_U17012_2;
    wire CHOR07_n_U17027_12;
    wire CHOR07_n_U24017_2;
    wire CHOR08_n;
    wire CHOR08_n_U16021_4;
    wire CHOR08_n_U17012_4;
    wire CHOR08_n_U17041_12;
    wire CHOR08_n_U24017_4;
    wire CHOR09_n;
    wire CHOR09_n_U17012_6;
    wire CHOR09_n_U17052_2;
    wire CHOR09_n_U24017_6;
    wire CHOR09_n_U24017_8;
    wire CHOR10_n;
    wire CHOR10_n_U17012_8;
    wire CHOR10_n_U17052_4;
    wire CHOR10_n_U24017_10;
    wire CHOR10_n_U24017_12;
    wire CHOR11_n;
    wire CHOR11_n_U17012_10;
    wire CHOR11_n_U17052_6;
    wire CHOR11_n_U24021_2;
    wire CHOR11_n_U24021_4;
    wire CHOR12_n;
    wire CHOR12_n_U17012_12;
    wire CHOR12_n_U17052_8;
    wire CHOR12_n_U24021_6;
    wire CHOR13_n;
    wire CHOR13_n_U17019_2;
    wire CHOR13_n_U17052_10;
    wire CHOR13_n_U24021_8;
    wire CHOR14_n;
    wire CHOR14_n_U17019_4;
    wire CHOR14_n_U17052_12;
    wire CHOR14_n_U24021_10;
    wire CHOR16_n;
    wire CHOR16_n_U17019_6;
    wire CHOR16_n_U17061_2;
    wire CHOR16_n_U24021_12;
    wire CHWL01_n;
    wire CHWL02_n;
    wire CHWL03_n;
    wire CHWL04_n;
    wire CHWL05_n;
    wire CHWL06_n;
    wire CHWL07_n;
    wire CHWL08_n;
    wire CHWL09_n;
    wire CHWL10_n;
    wire CHWL11_n;
    wire CHWL12_n;
    wire CHWL13_n;
    wire CHWL14_n;
    wire CHWL16_n;
    wire CI01_n;
    wire CI05_n;
    wire CI09_n;
    wire CI13_n;
    wire CI_n;
    wire CI_n_U4061_12;
    wire CI_n_U5018_2;
    wire CI_n_U5044_10;
    wire CI_n_U6047_2;
    wire CLG1G;
    wire CLG2G;
    wire CLROPE;
    wire CLXC;
    wire CO06;
    wire CO06_U8041_2;
    wire CO06_U8050_2;
    wire CO10;
    wire CO10_U9041_2;
    wire CO10_U9050_2;
    wire CO14;
    wire CO14_U10041_2;
    wire CO14_U10050_2;
    wire CQG;
    wire CSG;
    wire CT;
    wire CTROR;
    wire CTROR_n;
    wire CT_n;
    wire CUG;
    wire CXB0_n;
    wire CXB1_n;
    wire CXB2_n;
    wire CXB3_n;
    wire CXB4_n;
    wire CXB5_n;
    wire CXB6_n;
    wire CXB7_n;
    wire CYL_n;
    wire CYR_n;
    wire CZG;
    wire DAS0;
    wire DAS0_n;
    wire DAS1;
    wire DAS1_n;
    wire DCA0;
    wire DCS0;
    wire DIM0_n;
    wire DINC;
    wire DINC_n;
    wire DIVSTG;
    wire DIV_n;
    wire DLKPLS;
    wire DRPRST;
    wire DV1;
    wire DV1376;
    wire DV1376_n;
    wire DV1_n;
    wire DV3764;
    wire DV376_n;
    wire DV4;
    wire DV4B1B;
    wire DV4_n;
    wire DVST;
    wire DXCH0;
    wire E5;
    wire E6;
    wire E7_n;
    wire EAC_n;
    wire EB10;
    wire EB11_n;
    wire EB9;
    wire EDOP_n;
    wire EMSD;
    wire ERRST;
    wire EXST0_n;
    wire EXST1_n;
    wire EXT;
    wire EXTPLS;
    wire F01A;
    wire F01B;
    wire F02B;
    wire F03B;
    wire F04A;
    wire F04B;
    wire F05A_n;
    wire F05B_n;
    wire F06B;
    wire F07A;
    wire F07B;
    wire F07B_n;
    wire F08B;
    wire F09A;
    wire F09B;
    wire F09B_n;
    wire F10A;
    wire F10A_n;
    wire F10B;
    wire F12B;
    wire F14B;
    wire F17A;
    wire F17B;
    wire F18A;
    wire F18B;
    wire F5ASB0_n;
    wire F5ASB2;
    wire F5ASB2_n;
    wire F5BSB2_n;
    wire FETCH0;
    wire FETCH0_n;
    wire FETCH1;
    wire FLASH;
    wire FLASH_n;
    wire FS01;
    wire FS01_n;
    wire FS02;
    wire FS03;
    wire FS04;
    wire FS05;
    wire FS05_n;
    wire FS06;
    wire FS07A;
    wire FS07_n;
    wire FS08;
    wire FS09;
    wire FS09_n;
    wire FS10;
    wire FS13;
    wire FS14;
    wire FS16;
    wire FS17;
    wire FUTEXT;
    wire G01;
    wire G01ED;
    wire G01_n;
    wire G01_n_U8013_6;
    wire G01_n_U8013_8;
    wire G02;
    wire G02ED;
    wire G03;
    wire G03ED;
    wire G04;
    wire G04ED;
    wire G05;
    wire G05ED;
    wire G05_n;
    wire G05_n_U9013_6;
    wire G05_n_U9013_8;
    wire G06;
    wire G06ED;
    wire G06_n;
    wire G06_n_U9028_10;
    wire G06_n_U9028_12;
    wire G07;
    wire G07ED;
    wire G07_n;
    wire G07_n_U9050_6;
    wire G07_n_U9050_8;
    wire G08;
    wire G09;
    wire G09_n;
    wire G09_n_U10013_6;
    wire G09_n_U10013_8;
    wire G10;
    wire G10_n;
    wire G10_n_U10028_10;
    wire G10_n_U10028_12;
    wire G11;
    wire G11_n;
    wire G11_n_U10050_6;
    wire G11_n_U10050_8;
    wire G12;
    wire G13;
    wire G13_n;
    wire G13_n_U11013_6;
    wire G13_n_U11013_8;
    wire G14;
    wire G14_n;
    wire G14_n_U11028_10;
    wire G14_n_U11028_12;
    wire G15;
    wire G15_n;
    wire G15_n_U11050_6;
    wire G15_n_U11050_8;
    wire G16;
    wire G16SW_n;
    wire G2LSG_n;
    wire GEM01;
    wire GEM02;
    wire GEM03;
    wire GEM04;
    wire GEM05;
    wire GEM06;
    wire GEM07;
    wire GEM08;
    wire GEM09;
    wire GEM10;
    wire GEM11;
    wire GEM12;
    wire GEM13;
    wire GEM14;
    wire GEM16;
    wire GEMP;
    wire GEQZRO_n;
    wire GINH;
    wire GNHNC;
    wire GOJ1;
    wire GOJ1_n;
    wire GOJAM;
    wire GOJAM_n;
    wire GTONE;
    wire GTONE_U24029_2;
    wire GTONE_U24029_4;
    wire GTRST_n;
    wire GTSET;
    wire GTSET_n;
    wire GYROD;
    wire HIMOD;
    wire HNDRPT;
    wire IC1;
    wire IC10;
    wire IC10_n;
    wire IC11;
    wire IC11_n;
    wire IC12;
    wire IC12_n;
    wire IC13;
    wire IC14;
    wire IC15;
    wire IC15_n;
    wire IC16;
    wire IC16_n;
    wire IC17;
    wire IC2;
    wire IC2_n;
    wire IC3;
    wire IC4;
    wire IC5;
    wire IC5_n;
    wire IC6;
    wire IC7;
    wire IC8_n;
    wire IC9;
    wire IIP;
    wire IIP_n;
    wire IL01;
    wire IL02;
    wire IL03;
    wire IL04;
    wire IL05;
    wire IL06;
    wire IL07;
    wire INCR0;
    wire INCSET_n;
    wire INHPLS;
    wire INHPLS_U12016_10;
    wire INHPLS_U12016_12;
    wire INKL;
    wire INKL_n;
    wire INLNKM;
    wire INLNKP;
    wire INOTLD;
    wire INOUT;
    wire INOUT_n;
    wire KRPT;
    wire KYRPT1;
    wire KYRPT2;
    wire L01_n;
    wire L01_n_U8007_6;
    wire L02_n;
    wire L02_n_U8013_12;
    wire L04_n;
    wire L04_n_U8050_12;
    wire L08_n;
    wire L08_n_U9050_12;
    wire L12_n;
    wire L12_n_U10050_12;
    wire L15_n;
    wire L15_n_U11041_6;
    wire L16_n;
    wire L16_n_U11050_12;
    wire L16_n_U4063_8;
    wire L2GDG_n;
    wire L2GD_n;
    wire LOMOD;
    wire MASK0;
    wire MASK0_n;
    wire MBR1_U4066_8;
    wire MBR2_U4066_10;
    wire MCDU;
    wire MCRO_n;
    wire MCTRAL_n_U13051_12;
    wire MGOJAM_U2148_6;
    wire MIIP_U3053_6;
    wire MINC;
    wire MINHL_U3053_4;
    wire MINKL_U13053_4;
    wire MKRPT;
    wire MNISQ_U5068_2;
    wire MON800_U24038_2;
    wire MONEX;
    wire MONEX_n;
    wire MONEX_n_U5005_2;
    wire MONEX_n_U6029_6;
    wire MONWT_U2148_2;
    wire MON_n;
    wire MONpCH;
    wire MOSCAL_n_U13053_2;
    wire MOUT_n;
    wire MP0;
    wire MP0T10;
    wire MP0_n;
    wire MP1;
    wire MP1_n;
    wire MP3;
    wire MP3A;
    wire MP3_n;
    wire MPAL_n_U12050_2;
    wire MPIPAL_n_U13052_4;
    wire MRAG_U7040_2;
    wire MRCH_U6058_2;
    wire MREQIN_U13053_6;
    wire MRGG_U7039_12;
    wire MRLG_U7040_4;
    wire MRPTAL_n_U13051_8;
    wire MRSC_U4067_2;
    wire MRULOG_U7040_6;
    wire MSCAFL_n_U13052_10;
    wire MSCDBL_n_U13052_6;
    wire MSQ10_U3053_2;
    wire MSQ11_U3054_12;
    wire MSQ12_U3054_10;
    wire MSQ13_U3054_8;
    wire MSQ14_U3054_6;
    wire MSQ16_U3054_4;
    wire MSQEXT_U3054_2;
    wire MST1_U4066_2;
    wire MST2_U4066_4;
    wire MST3_U4066_6;
    wire MSTPIT_n_U2148_8;
    wire MSTRTP;
    wire MSU0;
    wire MSU0_n;
    wire MT01_U2046_2;
    wire MT02_U2046_4;
    wire MT03_U2046_6;
    wire MT04_U2046_8;
    wire MT05_U2046_10;
    wire MT06_U2046_12;
    wire MT07_U2047_2;
    wire MT08_U2047_4;
    wire MT09_U2047_6;
    wire MT10_U2047_8;
    wire MT11_U2047_10;
    wire MT12_U2047_12;
    wire MTCAL_n_U13051_10;
    wire MTCSA_n_U3053_8;
    wire MVFAIL_n_U13052_2;
    wire MWAG_U7038_12;
    wire MWARNF_n_U13052_12;
    wire MWATCH_n_U13052_8;
    wire MWBBEG_U7039_10;
    wire MWBG_U7038_4;
    wire MWCH_U4066_12;
    wire MWEBG_U7039_6;
    wire MWFBG_U7039_8;
    wire MWG_U7038_6;
    wire MWL01_U8068_2;
    wire MWL02_U8068_4;
    wire MWL03_U8068_6;
    wire MWL04_U8068_8;
    wire MWL05_U9068_2;
    wire MWL06_U9068_4;
    wire MWL07_U9068_6;
    wire MWL08_U9068_8;
    wire MWL09_U10068_2;
    wire MWL10_U10068_4;
    wire MWL11_U10068_6;
    wire MWL12_U10068_8;
    wire MWL13_U11068_2;
    wire MWL14_U11068_4;
    wire MWL15_U11068_6;
    wire MWL16_U11068_8;
    wire MWLG_U7038_10;
    wire MWQG_U7039_4;
    wire MWSG_U7039_2;
    wire MWYG_U7038_2;
    wire MWZG_U7038_8;
    wire NDR100_n;
    wire NDX0_n;
    wire NDXX1_n;
    wire NEAC;
    wire NISQ;
    wire NISQL_n;
    wire NISQ_n;
    wire OCTAD2;
    wire OCTAD3;
    wire OCTAD4;
    wire OCTAD5;
    wire OCTAD6;
    wire OSCALM;
    wire OTLNKM;
    wire OVF_n;
    wire P01;
    wire P01_n;
    wire P02;
    wire P02_n;
    wire P03;
    wire P03_n;
    wire P04;
    wire P04_n;
    wire P05;
    wire P05_n;
    wire PALE;
    wire PALE_U12027_2;
    wire PALE_U12027_4;
    wire PC15_n;
    wire PCDU;
    wire PHS2;
    wire PHS2_n;
    wire PHS3_n;
    wire PHS4;
    wire PHS4_n;
    wire PIFL_n;
    wire PINC;
    wire PIPAFL;
    wire PIPPLS_n;
    wire PIPXM;
    wire PIPXP;
    wire PIPYM;
    wire PIPYP;
    wire PIPZM;
    wire PIPZP;
    wire PONEX;
    wire POUT_n;
    wire PRINC;
    wire PSEUDO;
    wire PTWOX;
    wire QC0_n;
    wire QC1_n;
    wire QC2_n;
    wire QC3_n;
    wire QXCH0_n;
    wire R15;
    wire R1C;
    wire R1C_n;
    wire R1C_n_U4063_10;
    wire R1C_n_U6029_12;
    wire R6;
    wire RAD;
    wire RADRG;
    wire RADRPT;
    wire RADRZ;
    wire RAG_n;
    wire RAND0;
    wire RA_n;
    wire RA_n_U4039_10;
    wire RA_n_U4045_8;
    wire RA_n_U5005_8;
    wire RA_n_U5024_4;
    wire RA_n_U5039_12;
    wire RB1;
    wire RB1F;
    wire RB1_n;
    wire RB1_n_U4063_6;
    wire RB1_n_U6029_10;
    wire RB2;
    wire RBBEG_n;
    wire RBHG_n;
    wire RBLG_n;
    wire RBSQ;
    wire RB_n;
    wire RB_n_U4039_2;
    wire RB_n_U4061_10;
    wire RB_n_U5005_6;
    wire RB_n_U5018_10;
    wire RB_n_U5049_2;
    wire RB_n_U6004_8;
    wire RB_n_U6037_8;
    wire RCG_n;
    wire RCH11_n;
    wire RCH12_n;
    wire RCH13_n;
    wire RCH14_n;
    wire RCH33_n;
    wire RCHAT_n;
    wire RCHBT_n;
    wire RCHG_n;
    wire RCH_n;
    wire RC_n;
    wire RC_n_U4039_4;
    wire RC_n_U4061_8;
    wire RC_n_U5012_8;
    wire RC_n_U5024_10;
    wire RC_n_U5049_10;
    wire RC_n_U6047_6;
    wire RC_n_U6052_8;
    wire READ0;
    wire REBG_n;
    wire RELPLS;
    wire RELPLS_U12016_6;
    wire RELPLS_U12016_8;
    wire RESETA;
    wire RESETB;
    wire RESETC;
    wire RESETD;
    wire REX;
    wire REY;
    wire RFBG_n;
    wire RGG_n;
    wire RG_n;
    wire RG_n_U5012_6;
    wire RG_n_U5044_2;
    wire RG_n_U5044_4;
    wire RG_n_U5059_10;
    wire RG_n_U6014_8;
    wire RL01_n;
    wire RL01_n_U15039_12;
    wire RL01_n_U8007_10;
    wire RL01_n_U8007_12;
    wire RL01_n_U8007_4;
    wire RL01_n_U8013_4;
    wire RL02_n;
    wire RL02_n_U15039_10;
    wire RL02_n_U8013_10;
    wire RL02_n_U8028_2;
    wire RL02_n_U8028_6;
    wire RL02_n_U8028_8;
    wire RL03_n;
    wire RL03_n_U15039_4;
    wire RL03_n_U8041_10;
    wire RL03_n_U8041_12;
    wire RL03_n_U8041_4;
    wire RL03_n_U8050_4;
    wire RL04_n;
    wire RL04_n_U15039_6;
    wire RL04_n_U8050_10;
    wire RL04_n_U8061_2;
    wire RL04_n_U8061_6;
    wire RL04_n_U8061_8;
    wire RL05_n;
    wire RL05_n_U15039_8;
    wire RL05_n_U9007_10;
    wire RL05_n_U9007_12;
    wire RL05_n_U9007_4;
    wire RL05_n_U9013_4;
    wire RL06_n;
    wire RL06_n_U15016_6;
    wire RL06_n_U9013_10;
    wire RL06_n_U9028_2;
    wire RL06_n_U9028_6;
    wire RL06_n_U9028_8;
    wire RL09_n;
    wire RL09_n_U10007_10;
    wire RL09_n_U10007_12;
    wire RL09_n_U10007_4;
    wire RL09_n_U10013_4;
    wire RL09_n_U15016_4;
    wire RL10BB;
    wire RL10_n;
    wire RL10_n_U10013_10;
    wire RL10_n_U10028_2;
    wire RL10_n_U10028_6;
    wire RL10_n_U10028_8;
    wire RL10_n_U15016_2;
    wire RL11_n;
    wire RL11_n_U10041_10;
    wire RL11_n_U10041_12;
    wire RL11_n_U10041_4;
    wire RL11_n_U10050_4;
    wire RL11_n_U15004_12;
    wire RL12_n;
    wire RL12_n_U10050_10;
    wire RL12_n_U10061_2;
    wire RL12_n_U10061_6;
    wire RL12_n_U10061_8;
    wire RL12_n_U15004_10;
    wire RL13_n;
    wire RL13_n_U11007_10;
    wire RL13_n_U11007_12;
    wire RL13_n_U11007_4;
    wire RL13_n_U11013_4;
    wire RL13_n_U15004_8;
    wire RL14_n;
    wire RL14_n_U11013_10;
    wire RL14_n_U11028_2;
    wire RL14_n_U11028_6;
    wire RL14_n_U11028_8;
    wire RL14_n_U15004_6;
    wire RL15_n;
    wire RL15_n_U11041_10;
    wire RL15_n_U11041_12;
    wire RL15_n_U11041_4;
    wire RL15_n_U11050_4;
    wire RL15_n_U15004_4;
    wire RL16_n;
    wire RL16_n_U11050_10;
    wire RL16_n_U11061_2;
    wire RL16_n_U11061_6;
    wire RL16_n_U11061_8;
    wire RL16_n_U15004_2;
    wire RLG_n;
    wire RL_n;
    wire RL_n_U5005_12;
    wire RL_n_U5039_10;
    wire RNRADM;
    wire RNRADP;
    wire ROPER;
    wire ROPES;
    wire ROPET;
    wire ROR0;
    wire RPTSET;
    wire RPTSET_U3011_2;
    wire RPTSET_U3011_4;
    wire RPTSET_U3011_6;
    wire RPTSET_U6052_4;
    wire RQG_n;
    wire RQ_n;
    wire RRPA;
    wire RSCT;
    wire RSC_n;
    wire RSM3;
    wire RSM3_n;
    wire RSSB;
    wire RSTKX_n;
    wire RSTKY_n;
    wire RSTRT;
    wire RSTSTG;
    wire RT;
    wire RT_n;
    wire RUG_n;
    wire RULOG_n;
    wire RUPT0;
    wire RUPT1;
    wire RUPTOR_n;
    wire RUS_n;
    wire RU_n;
    wire RU_n_U5024_2;
    wire RU_n_U5059_4;
    wire RU_n_U5059_6;
    wire RU_n_U6014_12;
    wire RU_n_U6037_2;
    wire RU_n_U6052_6;
    wire RXOR0;
    wire RXOR0_n;
    wire RZG_n;
    wire RZ_n;
    wire RZ_n_U5005_4;
    wire RZ_n_U5018_4;
    wire RZ_n_U5049_4;
    wire RZ_n_U6052_2;
    wire S01;
    wire S01_n;
    wire S02;
    wire S02_n;
    wire S03;
    wire S03_n;
    wire S04;
    wire S04_n;
    wire S05;
    wire S05_n;
    wire S06;
    wire S06_n;
    wire S07;
    wire S07_n;
    wire S08;
    wire S08_n;
    wire S09;
    wire S09_n;
    wire S10;
    wire S10_n;
    wire S11;
    wire S11_n;
    wire S12;
    wire S12_n;
    wire SA01;
    wire SA01_U31001_29;
    wire SA01_U31023_16;
    wire SA01_U31025_7;
    wire SA02;
    wire SA02_U31001_31;
    wire SA02_U31023_14;
    wire SA02_U31025_8;
    wire SA03;
    wire SA03_U31001_33;
    wire SA03_U31023_12;
    wire SA03_U31025_9;
    wire SA04;
    wire SA04_U31001_35;
    wire SA04_U31023_9;
    wire SA04_U31025_10;
    wire SA05;
    wire SA05_U31001_38;
    wire SA05_U31023_7;
    wire SA05_U31025_13;
    wire SA06;
    wire SA06_U31001_40;
    wire SA06_U31023_5;
    wire SA06_U31025_14;
    wire SA07;
    wire SA07_U31001_42;
    wire SA07_U31023_3;
    wire SA07_U31025_15;
    wire SA08;
    wire SA08_U31001_44;
    wire SA08_U31024_18;
    wire SA08_U31025_16;
    wire SA09;
    wire SA09_U31001_30;
    wire SA09_U31024_16;
    wire SA09_U31025_29;
    wire SA10;
    wire SA10_U31001_32;
    wire SA10_U31024_14;
    wire SA10_U31025_30;
    wire SA11;
    wire SA11_U31001_34;
    wire SA11_U31024_12;
    wire SA11_U31025_31;
    wire SA12;
    wire SA12_U31001_36;
    wire SA12_U31024_9;
    wire SA12_U31025_32;
    wire SA13;
    wire SA13_U31001_39;
    wire SA13_U31024_7;
    wire SA13_U31025_35;
    wire SA14;
    wire SA14_U31001_41;
    wire SA14_U31024_5;
    wire SA14_U31025_36;
    wire SA16;
    wire SA16_U31001_45;
    wire SA16_U31024_3;
    wire SA16_U31025_38;
    wire SAP;
    wire SAP_U31001_43;
    wire SAP_U31023_18;
    wire SAP_U31025_37;
    wire SB0_n;
    wire SB1_n;
    wire SB2;
    wire SB2_n;
    wire SB4;
    wire SBE;
    wire SBF;
    wire SBY;
    wire SCAD;
    wire SCAD_U5049_6;
    wire SCAD_U5049_8;
    wire SCAD_n;
    wire SETAB;
    wire SETCD;
    wire SETEK;
    wire SHAFTD;
    wire SHANC_n;
    wire SHIFT;
    wire SHIFT_n;
    wire SHINC_n;
    wire SHFTDM;
    wire SHFTDP;
    wire SQ0_n;
    wire SQ1_n;
    wire SQ2_n;
    wire SQEXT;
    wire SQEXT_n;
    wire SQR10;
    wire SQR10_n;
    wire SQR12_n;
    wire SR_n;
    wire ST0_n;
    wire ST1;
    wire ST1_n;
    wire ST2;
    wire ST2_n;
    wire ST2_n_U5024_6;
    wire ST2_n_U6047_12;
    wire ST3_n;
    wire STBE;
    wire STBF;
    wire STD2;
    wire STFET1_n;
    wire STNDBY_n;
    wire STOP;
    wire STOPA;
    wire STOP_n;
    wire STORE1_n;
    wire STR14;
    wire STR19;
    wire STR210;
    wire STR311;
    wire STR412;
    wire STR58;
    wire STR912;
    wire STRGAT;
    wire STRT1;
    wire STRTFC;
    wire SU0;
    wire SUMA01_n;
    wire SUMA02_n;
    wire SUMA03_n;
    wire SUMA11_n;
    wire SUMA12_n;
    wire SUMA13_n;
    wire SUMA14_n;
    wire SUMA15_n;
    wire SUMA16_n;
    wire SUMB01_n;
    wire SUMB02_n;
    wire SUMB03_n;
    wire SUMB11_n;
    wire SUMB12_n;
    wire SUMB13_n;
    wire SUMB14_n;
    wire SUMB15_n;
    wire SUMB16_n;
    wire T01;
    wire T01_n;
    wire T02;
    wire T02_n;
    wire T03;
    wire T03_n;
    wire T04;
    wire T04_n;
    wire T05;
    wire T05_n;
    wire T06;
    wire T06_n;
    wire T07;
    wire T07_n;
    wire T08;
    wire T08_n;
    wire T09;
    wire T09_n;
    wire T10;
    wire T10_n;
    wire T11;
    wire T11_n;
    wire T12;
    wire T12A;
    wire T12USE_n;
    wire T12_n;
    wire T1P;
    wire T2P;
    wire T3P;
    wire T4P;
    wire T5P;
    wire T6ON_n;
    wire T6P;
    wire T6RPT;
    wire TC0;
    wire TC0_n;
    wire TCF0;
    wire TCSAJ3;
    wire TCSAJ3_n;
    wire THRSTD;
    wire TIMR;
    wire TL15;
    wire TMPOUT;
    wire TMZ_n;
    wire TMZ_n_U4045_12;
    wire TMZ_n_U5012_2;
    wire TMZ_n_U5065_6;
    wire TOV_n;
    wire TOV_n_U5059_2;
    wire TOV_n_U6019_4;
    wire TPARG_n;
    wire TPOR_n;
    wire TPZG_n;
    wire TRNDM;
    wire TRNDP;
    wire TRSM;
    wire TRUND;
    wire TS0;
    wire TS0_n;
    wire TSGN_n;
    wire TSGN_n_U4063_2;
    wire TSGN_n_U4063_4;
    wire TSGN_n_U5059_12;
    wire TSGN_n_U5065_10;
    wire TSGU_n;
    wire TSUDO_n;
    wire TT_n;
    wire TWOX;
    wire U2BBK;
    wire U2BBKG_n;
    wire UNF_n;
    wire UPRUPT;
    wire US2SG;
    wire WAG_n;
    wire WALSG_n;
    wire WAND0;
    wire WA_n;
    wire WA_n_U5005_10;
    wire WA_n_U5024_12;
    wire WA_n_U5056_6;
    wire WA_n_U6029_8;
    wire WA_n_U6047_4;
    wire WBBEG_n;
    wire WBG_n;
    wire WB_n;
    wire WB_n_U5018_12;
    wire WB_n_U5039_2;
    wire WB_n_U5039_4;
    wire WB_n_U5059_8;
    wire WB_n_U6014_10;
    wire WCH11_n;
    wire WCH12_n;
    wire WCH13_n;
    wire WCH14_n;
    wire WCH34_n;
    wire WCH35_n;
    wire WCHG_n;
    wire WCH_n;
    wire WEBG_n;
    wire WEDOPG_n;
    wire WEX;
    wire WEY;
    wire WFBG_n;
    wire WG1G_n;
    wire WG2G_n;
    wire WG3G_n;
    wire WG4G_n;
    wire WG5G_n;
    wire WG_n;
    wire WG_n_U4039_12;
    wire WG_n_U4045_10;
    wire WG_n_U4045_2;
    wire WG_n_U5012_4;
    wire WG_n_U6019_8;
    wire WG_n_U6037_6;
    wire WHOMP;
    wire WHOMPA;
    wire WL01;
    wire WL01_n;
    wire WL02;
    wire WL02_n;
    wire WL03;
    wire WL03_n;
    wire WL04;
    wire WL04_n;
    wire WL05;
    wire WL05_n;
    wire WL06;
    wire WL06_n;
    wire WL07;
    wire WL07_n;
    wire WL08;
    wire WL08_n;
    wire WL09;
    wire WL09_n;
    wire WL10;
    wire WL10_n;
    wire WL11;
    wire WL11_n;
    wire WL12;
    wire WL12_n;
    wire WL13;
    wire WL13_n;
    wire WL14;
    wire WL14_n;
    wire WL15;
    wire WL15_n;
    wire WL16;
    wire WL16_n;
    wire WLG_n;
    wire WL_n;
    wire WL_n_U4061_6;
    wire WL_n_U5065_4;
    wire WL_n_U6014_6;
    wire WOR0;
    wire WOVR_n;
    wire WQG_n;
    wire WQ_n;
    wire WSC_n;
    wire WSC_n_U6019_6;
    wire WSC_n_U6037_4;
    wire WSG_n;
    wire WS_n;
    wire WS_n_U5034_12;
    wire WS_n_U6041_8;
    wire WT;
    wire WT_n;
    wire WY12_n;
    wire WY12_n_U5018_6;
    wire WY12_n_U5044_12;
    wire WYDG_n;
    wire WYDLOG_n;
    wire WYD_n;
    wire WYD_n_U5065_8;
    wire WYD_n_U6004_10;
    wire WYHIG_n;
    wire WYLOG_n;
    wire WY_n;
    wire WY_n_U4061_2;
    wire WY_n_U4061_4;
    wire WY_n_U5012_12;
    wire WY_n_U5024_8;
    wire WY_n_U5044_6;
    wire WY_n_U6004_12;
    wire WZG_n;
    wire WZ_n;
    wire WZ_n_U5018_8;
    wire WZ_n_U5056_12;
    wire WZ_n_U6019_2;
    wire XB0;
    wire XB0_n;
    wire XB1;
    wire XB1E;
    wire XB1_n;
    wire XB2;
    wire XB2E;
    wire XB2_n;
    wire XB3;
    wire XB3E;
    wire XB3_n;
    wire XB4;
    wire XB4E;
    wire XB4_n;
    wire XB5;
    wire XB5E;
    wire XB5_n;
    wire XB6;
    wire XB6E;
    wire XB6_n;
    wire XB7;
    wire XB7E;
    wire XB7_n;
    wire XT0_n;
    wire XT1E;
    wire XT1_n;
    wire XT2E;
    wire XT2_n;
    wire XT3E;
    wire XT3_n;
    wire XT4E;
    wire XT4_n;
    wire XT5E;
    wire XT5_n;
    wire XT6E;
    wire XT6_n;
    wire XT7E;
    wire XUY01_n;
    wire XUY02_n;
    wire XUY05_n;
    wire XUY06_n;
    wire XUY09_n;
    wire XUY10_n;
    wire XUY13_n;
    wire XUY14_n;
    wire YB0_n;
    wire YB1E;
    wire YB2E;
    wire YB3E;
    wire YT0_n;
    wire YT1E;
    wire YT2E;
    wire YT3E;
    wire YT4E;
    wire YT5E;
    wire YT6E;
    wire YT7E;
    wire Z15_n;
    wire Z15_n_U11041_8;
    wire Z15_n_U5065_2;
    wire Z16_n;
    wire Z16_n_U11061_4;
    wire Z16_n_U5056_4;
    wire ZAP_n;
    wire ZID;
    wire ZOUT_n;
    wire __A01_1__F02A;
    wire __A01_1__F03A;
    wire __A01_1__F05A;
    wire __A01_1__F05B;
    wire __A01_1__F06A;
    wire __A01_1__F08A;
    wire __A01_1__F11A;
    wire __A01_1__F11B;
    wire __A01_1__F12A;
    wire __A01_1__F13A;
    wire __A01_1__F13B;
    wire __A01_1__F14A;
    wire __A01_1__F15A;
    wire __A01_1__F15B;
    wire __A01_1__F16A;
    wire __A01_1__F16B;
    wire __A01_1__FS02A;
    wire __A01_1__FS03A;
    wire __A01_1__FS04A;
    wire __A01_1__FS05A;
    wire __A01_1__FS07;
    wire __A01_1__FS11;
    wire __A01_1__FS12;
    wire __A01_1__FS15;
    wire __A01_1__scaler_s10__FS_n;
    wire __A01_1__scaler_s11__FS_n;
    wire __A01_1__scaler_s12__FS_n;
    wire __A01_1__scaler_s13__FS_n;
    wire __A01_1__scaler_s14__FS_n;
    wire __A01_1__scaler_s15__FS_n;
    wire __A01_1__scaler_s16__FS_n;
    wire __A01_1__scaler_s17__FS_n;
    wire __A01_1__scaler_s2__FS_n;
    wire __A01_1__scaler_s3__FS_n;
    wire __A01_1__scaler_s4__FS_n;
    wire __A01_1__scaler_s5__FS_n;
    wire __A01_1__scaler_s6__FS_n;
    wire __A01_1__scaler_s7__FS_n;
    wire __A01_1__scaler_s8__FS_n;
    wire __A01_1__scaler_s9__FS_n;
    wire __A01_2__F19A;
    wire __A01_2__F19B;
    wire __A01_2__F20A;
    wire __A01_2__F20B;
    wire __A01_2__F21A;
    wire __A01_2__F21B;
    wire __A01_2__F22A;
    wire __A01_2__F22B;
    wire __A01_2__F23A;
    wire __A01_2__F23B;
    wire __A01_2__F24A;
    wire __A01_2__F24B;
    wire __A01_2__F25A;
    wire __A01_2__F25B;
    wire __A01_2__F26A;
    wire __A01_2__F26B;
    wire __A01_2__F27A;
    wire __A01_2__F27B;
    wire __A01_2__F28A;
    wire __A01_2__F28B;
    wire __A01_2__F29A;
    wire __A01_2__F29B;
    wire __A01_2__F30A;
    wire __A01_2__F30B;
    wire __A01_2__F31A;
    wire __A01_2__F31B;
    wire __A01_2__F32A;
    wire __A01_2__F32B;
    wire __A01_2__F33A;
    wire __A01_2__F33B;
    wire __A01_2__FS18;
    wire __A01_2__FS19;
    wire __A01_2__FS20;
    wire __A01_2__FS21;
    wire __A01_2__FS22;
    wire __A01_2__FS23;
    wire __A01_2__FS24;
    wire __A01_2__FS25;
    wire __A01_2__FS26;
    wire __A01_2__FS27;
    wire __A01_2__FS28;
    wire __A01_2__FS29;
    wire __A01_2__FS30;
    wire __A01_2__FS31;
    wire __A01_2__FS32;
    wire __A01_2__FS33;
    wire __A01_2__scaler_s18__FS_n;
    wire __A01_2__scaler_s19__FS_n;
    wire __A01_2__scaler_s20__FS_n;
    wire __A01_2__scaler_s21__FS_n;
    wire __A01_2__scaler_s22__FS_n;
    wire __A01_2__scaler_s23__FS_n;
    wire __A01_2__scaler_s24__FS_n;
    wire __A01_2__scaler_s25__FS_n;
    wire __A01_2__scaler_s26__FS_n;
    wire __A01_2__scaler_s27__FS_n;
    wire __A01_2__scaler_s28__FS_n;
    wire __A01_2__scaler_s29__FS_n;
    wire __A01_2__scaler_s30__FS_n;
    wire __A01_2__scaler_s31__FS_n;
    wire __A01_2__scaler_s32__FS_n;
    wire __A01_2__scaler_s33__FS_n;
    wire __A01_NET_175;
    wire __A01_NET_176;
    wire __A01_NET_177;
    wire __A01_NET_178;
    wire __A01_NET_179;
    wire __A01_NET_180;
    wire __A01_NET_181;
    wire __A01_NET_182;
    wire __A01_NET_183;
    wire __A01_NET_184;
    wire __A01_NET_185;
    wire __A01_NET_186;
    wire __A01_NET_187;
    wire __A01_NET_188;
    wire __A01_NET_189;
    wire __A01_NET_190;
    wire __A01_NET_191;
    wire __A01_NET_192;
    wire __A01_NET_193;
    wire __A01_NET_194;
    wire __A01_NET_195;
    wire __A01_NET_196;
    wire __A01_NET_197;
    wire __A01_NET_198;
    wire __A01_NET_199;
    wire __A01_NET_200;
    wire __A01_NET_201;
    wire __A01_NET_202;
    wire __A01_NET_203;
    wire __A01_NET_204;
    wire __A01_NET_205;
    wire __A01_NET_206;
    wire __A01_NET_207;
    wire __A01_NET_208;
    wire __A01_NET_209;
    wire __A01_NET_210;
    wire __A01_NET_211;
    wire __A01_NET_212;
    wire __A01_NET_213;
    wire __A01_NET_214;
    wire __A01_NET_215;
    wire __A01_NET_216;
    wire __A01_NET_217;
    wire __A01_NET_218;
    wire __A01_NET_219;
    wire __A01_NET_220;
    wire __A01_NET_221;
    wire __A01_NET_222;
    wire __A01_NET_223;
    wire __A01_NET_224;
    wire __A01_NET_225;
    wire __A01_NET_226;
    wire __A01_NET_227;
    wire __A01_NET_228;
    wire __A01_NET_229;
    wire __A01_NET_230;
    wire __A01_NET_231;
    wire __A01_NET_232;
    wire __A01_NET_233;
    wire __A01_NET_234;
    wire __A01_NET_235;
    wire __A01_NET_236;
    wire __A01_NET_237;
    wire __A01_NET_238;
    wire __A02_1__EVNSET_n;
    wire __A02_1__ODDSET_n;
    wire __A02_1__OVFSTB_n;
    wire __A02_1__Q2A;
    wire __A02_1__Q2A_U2148_4;
    wire __A02_1__RINGA_n;
    wire __A02_1__RINGB_n;
    wire __A02_1__cdiv_1__A;
    wire __A02_1__cdiv_1__B;
    wire __A02_1__cdiv_1__D;
    wire __A02_1__cdiv_1__FS;
    wire __A02_1__cdiv_1__FS_n;
    wire __A02_1__cdiv_2__A;
    wire __A02_1__cdiv_2__B;
    wire __A02_1__cdiv_2__C;
    wire __A02_1__cdiv_2__D;
    wire __A02_1__cdiv_2__F;
    wire __A02_1__cdiv_2__FS;
    wire __A02_1__cdiv_2__FS_n;
    wire __A02_1__evnset;
    wire __A02_1__oddset;
    wire __A02_1__ovfstb_r1;
    wire __A02_1__ovfstb_r2;
    wire __A02_1__ovfstb_r3;
    wire __A02_1__ovfstb_r4;
    wire __A02_1__ovfstb_r5;
    wire __A02_1__ovfstb_r6;
    wire __A02_2__EDSET;
    wire __A02_2__F01C;
    wire __A02_2__F01D;
    wire __A02_2__SB0;
    wire __A02_2__SB1;
    wire __A02_2__T12DC_n;
    wire __A02_3__OVF;
    wire __A02_3__T01DC_n;
    wire __A02_3__T02DC_n;
    wire __A02_3__T03DC_n;
    wire __A02_3__T04DC_n;
    wire __A02_3__T05DC_n;
    wire __A02_3__T06DC_n;
    wire __A02_3__T07DC_n;
    wire __A02_3__T08DC_n;
    wire __A02_3__T09DC_n;
    wire __A02_3__T10DC_n;
    wire __A02_3__T12SET;
    wire __A02_3__T12SET_U2038_2;
    wire __A02_3__T12SET_U2038_4;
    wire __A02_3__T12SET_U2038_6;
    wire __A02_3__T12SET_U2038_8;
    wire __A02_3__UNF;
    wire __A02_NET_133;
    wire __A02_NET_142;
    wire __A02_NET_143;
    wire __A02_NET_144;
    wire __A02_NET_145;
    wire __A02_NET_146;
    wire __A02_NET_147;
    wire __A02_NET_148;
    wire __A02_NET_149;
    wire __A02_NET_150;
    wire __A02_NET_151;
    wire __A02_NET_151_U2120_2;
    wire __A02_NET_151_U2120_4;
    wire __A02_NET_152;
    wire __A02_NET_153;
    wire __A02_NET_154;
    wire __A02_NET_156;
    wire __A02_NET_158;
    wire __A02_NET_159;
    wire __A02_NET_160;
    wire __A02_NET_161;
    wire __A02_NET_162;
    wire __A02_NET_163;
    wire __A02_NET_164;
    wire __A02_NET_165;
    wire __A02_NET_166;
    wire __A02_NET_167;
    wire __A02_NET_168;
    wire __A02_NET_169;
    wire __A02_NET_170;
    wire __A02_NET_171;
    wire __A02_NET_172;
    wire __A02_NET_173;
    wire __A02_NET_174;
    wire __A02_NET_175;
    wire __A02_NET_176;
    wire __A02_NET_177;
    wire __A02_NET_178;
    wire __A02_NET_179;
    wire __A02_NET_180;
    wire __A02_NET_181;
    wire __A02_NET_182;
    wire __A02_NET_183;
    wire __A02_NET_184;
    wire __A02_NET_185;
    wire __A02_NET_186;
    wire __A02_NET_187;
    wire __A02_NET_188;
    wire __A02_NET_189;
    wire __A02_NET_190;
    wire __A02_NET_191;
    wire __A02_NET_192;
    wire __A02_NET_193;
    wire __A02_NET_194;
    wire __A02_NET_195;
    wire __A02_NET_196;
    wire __A02_NET_197;
    wire __A02_NET_198;
    wire __A02_NET_199;
    wire __A03_1__CSQG;
    wire __A03_1__INHINT;
    wire __A03_1__INKBT1;
    wire __A03_1__NISQL;
    wire __A03_1__OVNHRP;
    wire __A03_1__QC0;
    wire __A03_1__RPTFRC;
    wire __A03_1__SQ3_n;
    wire __A03_1__SQ4_n;
    wire __A03_1__SQ5_n;
    wire __A03_1__SQ6_n;
    wire __A03_1__SQ7_n;
    wire __A03_1__SQR11;
    wire __A03_1__SQR12;
    wire __A03_1__SQR13;
    wire __A03_1__SQR14;
    wire __A03_1__SQR16;
    wire __A03_1__WSQG_n;
    wire __A03_1__wsqg;
    wire __A03_2__AUG0;
    wire __A03_2__BMF0;
    wire __A03_2__BMF0_n;
    wire __A03_2__BZF0;
    wire __A03_2__BZF0_n;
    wire __A03_2__DIM0;
    wire __A03_2__IC13_n;
    wire __A03_2__IC13_n_U3011_10;
    wire __A03_2__IC13_n_U3011_8;
    wire __A03_2__IC3_n;
    wire __A03_2__IC4_n;
    wire __A03_2__IC9_n;
    wire __A03_2__LXCH0;
    wire __A03_2__NDX0;
    wire __A03_2__NDXX1;
    wire __A03_2__NEXST0;
    wire __A03_2__NEXST0_n;
    wire __A03_2__QXCH0;
    wire __A03_2__SQ5QC0_n;
    wire __A03_NET_163;
    wire __A03_NET_164;
    wire __A03_NET_165;
    wire __A03_NET_166;
    wire __A03_NET_167;
    wire __A03_NET_168;
    wire __A03_NET_169;
    wire __A03_NET_170;
    wire __A03_NET_171;
    wire __A03_NET_172;
    wire __A03_NET_173;
    wire __A03_NET_174;
    wire __A03_NET_175;
    wire __A03_NET_176;
    wire __A03_NET_177;
    wire __A03_NET_178;
    wire __A03_NET_179;
    wire __A03_NET_180;
    wire __A03_NET_181;
    wire __A03_NET_182;
    wire __A03_NET_183;
    wire __A03_NET_184;
    wire __A03_NET_185;
    wire __A03_NET_186;
    wire __A03_NET_187;
    wire __A03_NET_188;
    wire __A03_NET_189;
    wire __A03_NET_190;
    wire __A03_NET_191;
    wire __A03_NET_192;
    wire __A03_NET_193;
    wire __A03_NET_194;
    wire __A03_NET_196;
    wire __A03_NET_197;
    wire __A03_NET_198;
    wire __A03_NET_199;
    wire __A03_NET_200;
    wire __A03_NET_201;
    wire __A03_NET_202;
    wire __A03_NET_203;
    wire __A03_NET_204;
    wire __A03_NET_205;
    wire __A03_NET_206;
    wire __A03_NET_207;
    wire __A03_NET_208;
    wire __A03_NET_209;
    wire __A03_NET_211;
    wire __A03_NET_213;
    wire __A03_NET_214;
    wire __A03_NET_215;
    wire __A03_NET_216;
    wire __A03_NET_217;
    wire __A03_NET_218;
    wire __A03_NET_219;
    wire __A03_NET_220;
    wire __A03_NET_221;
    wire __A03_NET_223;
    wire __A03_NET_224;
    wire __A03_NET_225;
    wire __A03_NET_226;
    wire __A03_NET_227;
    wire __A03_NET_228;
    wire __A03_NET_231;
    wire __A03_NET_232;
    wire __A03_NET_234;
    wire __A03_NET_235;
    wire __A03_NET_236;
    wire __A03_NET_237;
    wire __A03_NET_238;
    wire __A03_NET_239;
    wire __A03_NET_240;
    wire __A03_NET_242;
    wire __A04_1__DV0;
    wire __A04_1__DV0_n;
    wire __A04_1__DV376;
    wire __A04_1__DVST_n;
    wire __A04_1__SGUM;
    wire __A04_1__SGUM_U4003_10;
    wire __A04_1__SGUM_U4003_12;
    wire __A04_1__ST1376_n;
    wire __A04_1__ST376;
    wire __A04_1__ST376_n;
    wire __A04_1__ST4_n;
    wire __A04_1__STG1;
    wire __A04_1__STG2;
    wire __A04_1__STG3;
    wire __A04_1__TRSM_n;
    wire __A04_1__TSGN2;
    wire __A04_2__BR12B;
    wire __A04_2__BR1B2;
    wire __A04_2__BRXP3;
    wire __A04_2__READ0_n;
    wire __A04_2__RUPT0_n;
    wire __A04_2__RUPT1_n;
    wire __A04_2__WOR0_n;
    wire __A04_2__WRITE0;
    wire __A04_2__WRITE0_n;
    wire __A04_NET_184;
    wire __A04_NET_185;
    wire __A04_NET_186;
    wire __A04_NET_187;
    wire __A04_NET_188;
    wire __A04_NET_189;
    wire __A04_NET_192;
    wire __A04_NET_193;
    wire __A04_NET_193_U4023_6;
    wire __A04_NET_193_U4023_8;
    wire __A04_NET_194;
    wire __A04_NET_195;
    wire __A04_NET_196;
    wire __A04_NET_197;
    wire __A04_NET_198;
    wire __A04_NET_199;
    wire __A04_NET_200;
    wire __A04_NET_201;
    wire __A04_NET_202;
    wire __A04_NET_203;
    wire __A04_NET_204;
    wire __A04_NET_204_U4023_10;
    wire __A04_NET_204_U4023_12;
    wire __A04_NET_204_U4029_2;
    wire __A04_NET_204_U4029_4;
    wire __A04_NET_204_U4029_6;
    wire __A04_NET_205;
    wire __A04_NET_206;
    wire __A04_NET_207;
    wire __A04_NET_208;
    wire __A04_NET_208_U4029_10;
    wire __A04_NET_208_U4029_8;
    wire __A04_NET_209;
    wire __A04_NET_210;
    wire __A04_NET_211;
    wire __A04_NET_214;
    wire __A04_NET_215;
    wire __A04_NET_215_U4023_2;
    wire __A04_NET_215_U4023_4;
    wire __A04_NET_222;
    wire __A04_NET_223;
    wire __A04_NET_225;
    wire __A04_NET_226;
    wire __A04_NET_227;
    wire __A04_NET_230;
    wire __A04_NET_231;
    wire __A04_NET_232;
    wire __A04_NET_233;
    wire __A04_NET_234;
    wire __A04_NET_235;
    wire __A04_NET_236;
    wire __A04_NET_236_U4003_6;
    wire __A04_NET_236_U4003_8;
    wire __A04_NET_237;
    wire __A04_NET_238;
    wire __A04_NET_239;
    wire __A04_NET_241;
    wire __A04_NET_244;
    wire __A04_NET_245;
    wire __A04_NET_246;
    wire __A04_NET_247;
    wire __A04_NET_248;
    wire __A04_NET_249;
    wire __A04_NET_249_U4003_2;
    wire __A04_NET_249_U4003_4;
    wire __A04_NET_250;
    wire __A04_NET_251;
    wire __A04_NET_252;
    wire __A04_NET_253;
    wire __A04_NET_254;
    wire __A04_NET_255;
    wire __A04_NET_256;
    wire __A04_NET_257;
    wire __A04_NET_258;
    wire __A04_NET_259;
    wire __A04_NET_260;
    wire __A04_NET_261;
    wire __A04_NET_262;
    wire __A04_NET_263;
    wire __A04_NET_266;
    wire __A04_NET_269;
    wire __A04_NET_270;
    wire __A04_NET_271;
    wire __A04_NET_272;
    wire __A04_NET_273;
    wire __A04_NET_274;
    wire __A04_NET_275;
    wire __A04_NET_276;
    wire __A04_NET_277;
    wire __A04_NET_278;
    wire __A04_NET_279;
    wire __A04_NET_279_U4045_4;
    wire __A04_NET_279_U4045_6;
    wire __A04_NET_280;
    wire __A04_NET_281;
    wire __A04_NET_282;
    wire __A04_NET_283;
    wire __A04_NET_284;
    wire __A04_NET_285;
    wire __A04_NET_286;
    wire __A04_NET_287;
    wire __A04_NET_288;
    wire __A04_NET_289;
    wire __A04_NET_290;
    wire __A04_NET_291;
    wire __A04_NET_292;
    wire __A04_NET_293;
    wire __A04_NET_294;
    wire __A04_NET_295;
    wire __A04_NET_296;
    wire __A04_NET_297;
    wire __A04_NET_298;
    wire __A04_NET_299;
    wire __A04_NET_300;
    wire __A04_NET_301;
    wire __A04_NET_302;
    wire __A04_NET_303;
    wire __A04_NET_304;
    wire __A04_NET_305;
    wire __A04_NET_306;
    wire __A04_NET_307;
    wire __A04_NET_308;
    wire __A04_NET_309;
    wire __A04_NET_310;
    wire __A04_NET_311;
    wire __A04_NET_312;
    wire __A04_NET_313;
    wire __A04_NET_314;
    wire __A04_NET_315;
    wire __A04_NET_316;
    wire __A04_NET_319;
    wire __A04_NET_320;
    wire __A04_NET_321;
    wire __A04_NET_322;
    wire __A04_NET_323;
    wire __A04_NET_324;
    wire __A04_NET_325;
    wire __A04_NET_326;
    wire __A04_NET_327;
    wire __A04_NET_328;
    wire __A04_NET_329;
    wire __A04_NET_334;
    wire __A04_NET_335;
    wire __A04_NET_336;
    wire __A04_NET_337;
    wire __A05_1__10XP6;
    wire __A05_1__10XP7;
    wire __A05_1__3XP5;
    wire __A05_1__8XP12;
    wire __A05_1__8XP15;
    wire __A05_1__8XP3;
    wire __A05_1__DV1B1B;
    wire __A05_1__PARTC;
    wire __A05_2__10XP10;
    wire __A05_2__11XP6;
    wire __A05_2__5XP13;
    wire __A05_2__5XP19;
    wire __A05_2__5XP9;
    wire __A05_2__6XP2;
    wire __A05_2__6XP7;
    wire __A05_NET_177;
    wire __A05_NET_178;
    wire __A05_NET_179;
    wire __A05_NET_181;
    wire __A05_NET_182;
    wire __A05_NET_183;
    wire __A05_NET_184;
    wire __A05_NET_185;
    wire __A05_NET_186;
    wire __A05_NET_187;
    wire __A05_NET_188;
    wire __A05_NET_189;
    wire __A05_NET_190;
    wire __A05_NET_191;
    wire __A05_NET_192;
    wire __A05_NET_193;
    wire __A05_NET_194;
    wire __A05_NET_196;
    wire __A05_NET_198;
    wire __A05_NET_199;
    wire __A05_NET_203;
    wire __A05_NET_204;
    wire __A05_NET_205;
    wire __A05_NET_206;
    wire __A05_NET_208;
    wire __A05_NET_209;
    wire __A05_NET_210;
    wire __A05_NET_211;
    wire __A05_NET_212;
    wire __A05_NET_213;
    wire __A05_NET_214;
    wire __A05_NET_215;
    wire __A05_NET_216;
    wire __A05_NET_217;
    wire __A05_NET_218;
    wire __A05_NET_219;
    wire __A05_NET_220;
    wire __A05_NET_221;
    wire __A05_NET_222;
    wire __A05_NET_223;
    wire __A05_NET_224;
    wire __A05_NET_225;
    wire __A05_NET_226;
    wire __A05_NET_227;
    wire __A05_NET_228;
    wire __A05_NET_229;
    wire __A05_NET_230;
    wire __A05_NET_231;
    wire __A05_NET_232;
    wire __A05_NET_233;
    wire __A05_NET_234;
    wire __A05_NET_235;
    wire __A05_NET_236;
    wire __A05_NET_237;
    wire __A05_NET_238;
    wire __A05_NET_239;
    wire __A05_NET_240;
    wire __A05_NET_243;
    wire __A05_NET_244;
    wire __A05_NET_245;
    wire __A05_NET_246;
    wire __A05_NET_247;
    wire __A05_NET_248;
    wire __A05_NET_249;
    wire __A05_NET_250;
    wire __A05_NET_251;
    wire __A05_NET_252;
    wire __A05_NET_253;
    wire __A05_NET_254;
    wire __A05_NET_255;
    wire __A05_NET_256;
    wire __A05_NET_257;
    wire __A05_NET_258;
    wire __A05_NET_259;
    wire __A05_NET_260;
    wire __A05_NET_260_U5049_12;
    wire __A05_NET_260_U5056_2;
    wire __A05_NET_261;
    wire __A05_NET_262;
    wire __A05_NET_263;
    wire __A05_NET_264;
    wire __A05_NET_265;
    wire __A05_NET_266;
    wire __A05_NET_267;
    wire __A05_NET_267_U5056_10;
    wire __A05_NET_267_U5056_8;
    wire __A05_NET_268;
    wire __A05_NET_269;
    wire __A05_NET_270;
    wire __A05_NET_271;
    wire __A05_NET_272;
    wire __A05_NET_273;
    wire __A05_NET_276;
    wire __A05_NET_277;
    wire __A05_NET_279;
    wire __A05_NET_280;
    wire __A05_NET_281;
    wire __A05_NET_282;
    wire __A05_NET_282_U5034_10;
    wire __A05_NET_282_U5034_8;
    wire __A05_NET_283;
    wire __A05_NET_284;
    wire __A05_NET_285;
    wire __A05_NET_285_U5039_6;
    wire __A05_NET_285_U5039_8;
    wire __A05_NET_286;
    wire __A05_NET_287;
    wire __A05_NET_288;
    wire __A05_NET_289;
    wire __A05_NET_291;
    wire __A05_NET_292;
    wire __A05_NET_293;
    wire __A05_NET_294;
    wire __A05_NET_296;
    wire __A05_NET_297;
    wire __A05_NET_298;
    wire __A05_NET_299;
    wire __A05_NET_300;
    wire __A05_NET_301;
    wire __A05_NET_302;
    wire __A05_NET_303;
    wire __A05_NET_305;
    wire __A05_NET_306;
    wire __A05_NET_307;
    wire __A05_NET_308;
    wire __A05_NET_309;
    wire __A05_NET_310;
    wire __A05_NET_313;
    wire __A05_NET_314;
    wire __A05_NET_315;
    wire __A05_NET_316;
    wire __A05_NET_317;
    wire __A05_NET_318;
    wire __A05_NET_319;
    wire __A05_NET_320;
    wire __A05_NET_323;
    wire __A05_NET_324;
    wire __A05_NET_325;
    wire __A05_NET_326;
    wire __A05_NET_327;
    wire __A05_NET_328;
    wire __A05_NET_330;
    wire __A05_NET_331;
    wire __A05_NET_333;
    wire __A05_NET_334;
    wire __A05_NET_335;
    wire __A05_NET_338;
    wire __A05_NET_339;
    wire __A05_NET_340;
    wire __A05_NET_341;
    wire __A05_NET_342;
    wire __A05_NET_343;
    wire __A05_NET_344;
    wire __A05_NET_345;
    wire __A05_NET_346;
    wire __A05_NET_348;
    wire __A05_NET_349;
    wire __A05_NET_350;
    wire __A05_NET_351;
    wire __A05_NET_352;
    wire __A06_1__DVXP1;
    wire __A06_1__L02A_n;
    wire __A06_1__WHOMP_n;
    wire __A06_1__ZAP;
    wire __A06_1__ZIP;
    wire __A06_1__ZIPCI;
    wire __A06_2__10XP15;
    wire __A06_2__10XP9;
    wire __A06_2__6XP10;
    wire __A06_2__6XP12;
    wire __A06_2__7XP10;
    wire __A06_2__7XP11;
    wire __A06_2__7XP15;
    wire __A06_2__7XP7;
    wire __A06_2__8XP4;
    wire __A06_2__MOUT;
    wire __A06_2__POUT;
    wire __A06_2__RDBANK;
    wire __A06_2__ZOUT;
    wire __A06_NET_183;
    wire __A06_NET_184;
    wire __A06_NET_185;
    wire __A06_NET_186;
    wire __A06_NET_186_U6041_10;
    wire __A06_NET_186_U6041_12;
    wire __A06_NET_190;
    wire __A06_NET_191;
    wire __A06_NET_192;
    wire __A06_NET_193;
    wire __A06_NET_195;
    wire __A06_NET_196;
    wire __A06_NET_197;
    wire __A06_NET_198;
    wire __A06_NET_199;
    wire __A06_NET_199_U6041_4;
    wire __A06_NET_199_U6041_6;
    wire __A06_NET_200;
    wire __A06_NET_203;
    wire __A06_NET_203_U6019_10;
    wire __A06_NET_203_U6019_12;
    wire __A06_NET_204;
    wire __A06_NET_205;
    wire __A06_NET_206;
    wire __A06_NET_207;
    wire __A06_NET_208;
    wire __A06_NET_209;
    wire __A06_NET_210;
    wire __A06_NET_211;
    wire __A06_NET_213;
    wire __A06_NET_214;
    wire __A06_NET_215;
    wire __A06_NET_216;
    wire __A06_NET_217;
    wire __A06_NET_219;
    wire __A06_NET_220;
    wire __A06_NET_220_U6047_10;
    wire __A06_NET_220_U6047_8;
    wire __A06_NET_221;
    wire __A06_NET_222;
    wire __A06_NET_223;
    wire __A06_NET_224;
    wire __A06_NET_226;
    wire __A06_NET_228;
    wire __A06_NET_229;
    wire __A06_NET_230;
    wire __A06_NET_231;
    wire __A06_NET_232;
    wire __A06_NET_233;
    wire __A06_NET_234;
    wire __A06_NET_236;
    wire __A06_NET_239;
    wire __A06_NET_240;
    wire __A06_NET_241;
    wire __A06_NET_241_U6029_2;
    wire __A06_NET_241_U6029_4;
    wire __A06_NET_242;
    wire __A06_NET_243;
    wire __A06_NET_244;
    wire __A06_NET_245;
    wire __A06_NET_246;
    wire __A06_NET_247;
    wire __A06_NET_248;
    wire __A06_NET_249;
    wire __A06_NET_250;
    wire __A06_NET_251;
    wire __A06_NET_253;
    wire __A06_NET_255;
    wire __A06_NET_256;
    wire __A06_NET_257;
    wire __A06_NET_258;
    wire __A06_NET_262;
    wire __A06_NET_264;
    wire __A06_NET_265;
    wire __A06_NET_266;
    wire __A06_NET_267;
    wire __A06_NET_268;
    wire __A06_NET_269;
    wire __A06_NET_270;
    wire __A06_NET_271;
    wire __A06_NET_272;
    wire __A06_NET_272_U6004_2;
    wire __A06_NET_272_U6004_4;
    wire __A06_NET_273;
    wire __A06_NET_274;
    wire __A06_NET_275;
    wire __A06_NET_276;
    wire __A06_NET_277;
    wire __A06_NET_280;
    wire __A06_NET_283;
    wire __A06_NET_284;
    wire __A06_NET_287;
    wire __A06_NET_288;
    wire __A06_NET_289;
    wire __A06_NET_290;
    wire __A06_NET_291;
    wire __A06_NET_292;
    wire __A06_NET_293;
    wire __A06_NET_294;
    wire __A06_NET_295;
    wire __A06_NET_296;
    wire __A06_NET_297;
    wire __A06_NET_298;
    wire __A06_NET_299;
    wire __A06_NET_300;
    wire __A06_NET_301;
    wire __A06_NET_302;
    wire __A06_NET_303;
    wire __A06_NET_304;
    wire __A06_NET_305;
    wire __A06_NET_306;
    wire __A06_NET_307;
    wire __A06_NET_308;
    wire __A06_NET_309;
    wire __A06_NET_310;
    wire __A06_NET_311;
    wire __A06_NET_312;
    wire __A06_NET_313;
    wire __A06_NET_314;
    wire __A06_NET_315;
    wire __A06_NET_316;
    wire __A06_NET_317;
    wire __A06_NET_318;
    wire __A06_NET_319;
    wire __A06_NET_320;
    wire __A06_NET_320_U6014_2;
    wire __A06_NET_320_U6014_4;
    wire __A06_NET_321;
    wire __A06_NET_322;
    wire __A06_NET_323;
    wire __A06_NET_324;
    wire __A06_NET_325;
    wire __A06_NET_326;
    wire __A06_NET_327;
    wire __A06_NET_328;
    wire __A06_NET_329;
    wire __A06_NET_330;
    wire __A06_NET_331;
    wire __A06_NET_332;
    wire __A06_NET_333;
    wire __A06_NET_334;
    wire __A06_NET_335;
    wire __A06_NET_336;
    wire __A06_NET_337;
    wire __A06_NET_339;
    wire __A06_NET_341;
    wire __A06_NET_345;
    wire __A06_NET_346;
    wire __A06_NET_347;
    wire __A06_NET_348;
    wire __A06_NET_350;
    wire __A06_NET_351;
    wire __A06_NET_352;
    wire __A07_1__WALSG;
    wire __A07_1__WGA_n;
    wire __A07_1__WGNORM;
    wire __A07_1__WSCG_n;
    wire __A07_2__CIFF;
    wire __A07_2__CINORM;
    wire __A07_2__G2LSG;
    wire __A07_2__RBBK;
    wire __A07_2__RSCG_n;
    wire __A07_2__RUSG_n;
    wire __A07_NET_133;
    wire __A07_NET_134;
    wire __A07_NET_135;
    wire __A07_NET_136;
    wire __A07_NET_137;
    wire __A07_NET_138;
    wire __A07_NET_139;
    wire __A07_NET_140;
    wire __A07_NET_143;
    wire __A07_NET_146;
    wire __A07_NET_147;
    wire __A07_NET_148;
    wire __A07_NET_149;
    wire __A07_NET_150;
    wire __A07_NET_151;
    wire __A07_NET_152;
    wire __A07_NET_153;
    wire __A07_NET_154;
    wire __A07_NET_155;
    wire __A07_NET_156;
    wire __A07_NET_157;
    wire __A07_NET_158;
    wire __A07_NET_158_U7007_2;
    wire __A07_NET_158_U7007_4;
    wire __A07_NET_159;
    wire __A07_NET_160;
    wire __A07_NET_161;
    wire __A07_NET_162;
    wire __A07_NET_163;
    wire __A07_NET_164;
    wire __A07_NET_165;
    wire __A07_NET_166;
    wire __A07_NET_167;
    wire __A07_NET_168;
    wire __A07_NET_170;
    wire __A07_NET_171;
    wire __A07_NET_172;
    wire __A07_NET_173;
    wire __A07_NET_174;
    wire __A07_NET_176;
    wire __A07_NET_177;
    wire __A07_NET_178;
    wire __A07_NET_179;
    wire __A07_NET_180;
    wire __A07_NET_181;
    wire __A07_NET_182;
    wire __A07_NET_183;
    wire __A07_NET_184;
    wire __A07_NET_186;
    wire __A07_NET_187;
    wire __A07_NET_188;
    wire __A07_NET_189;
    wire __A07_NET_190;
    wire __A07_NET_191;
    wire __A07_NET_194;
    wire __A07_NET_195;
    wire __A07_NET_196;
    wire __A07_NET_197;
    wire __A07_NET_198;
    wire __A07_NET_199;
    wire __A07_NET_200;
    wire __A07_NET_201;
    wire __A07_NET_202;
    wire __A07_NET_203;
    wire __A07_NET_204;
    wire __A07_NET_206;
    wire __A07_NET_207;
    wire __A07_NET_208;
    wire __A07_NET_209;
    wire __A07_NET_210;
    wire __A08_1__X1;
    wire __A08_1__X1_n;
    wire __A08_1__X2;
    wire __A08_1__X2_n;
    wire __A08_1__Y1;
    wire __A08_1__Y1_n;
    wire __A08_1__Y2;
    wire __A08_1__Y2_n;
    wire __A08_1___A1_n;
    wire __A08_1___A2_n;
    wire __A08_1___B1_n;
    wire __A08_1___B2_n;
    wire __A08_1___CI_INTERNAL;
    wire __A08_1___G2_n;
    wire __A08_1___G2_n_U8028_10;
    wire __A08_1___G2_n_U8028_12;
    wire __A08_1___Q1_n;
    wire __A08_1___Q2_n;
    wire __A08_1___RL_OUT_1;
    wire __A08_1___RL_OUT_2;
    wire __A08_1___Z1_n;
    wire __A08_1___Z1_n_U8007_8;
    wire __A08_1___Z2_n;
    wire __A08_1___Z2_n_U8028_4;
    wire __A08_2__X1;
    wire __A08_2__X1_n;
    wire __A08_2__X2;
    wire __A08_2__X2_n;
    wire __A08_2__Y1;
    wire __A08_2__Y1_n;
    wire __A08_2__Y2;
    wire __A08_2__Y2_n;
    wire __A08_2___A1_n;
    wire __A08_2___A2_n;
    wire __A08_2___B1_n;
    wire __A08_2___B2_n;
    wire __A08_2___CI_INTERNAL;
    wire __A08_2___G1_n;
    wire __A08_2___G1_n_U8050_6;
    wire __A08_2___G1_n_U8050_8;
    wire __A08_2___Q1_n;
    wire __A08_2___Q2_n;
    wire __A08_2___RL_OUT_1;
    wire __A08_2___RL_OUT_2;
    wire __A08_2___SUMA2;
    wire __A08_2___SUMB2;
    wire __A08_2___Z1_n;
    wire __A08_2___Z1_n_U8041_8;
    wire __A08_2___Z2_n;
    wire __A08_2___Z2_n_U8061_4;
    wire __A08_NET_137;
    wire __A08_NET_138;
    wire __A08_NET_139;
    wire __A08_NET_140;
    wire __A08_NET_141;
    wire __A08_NET_142;
    wire __A08_NET_143;
    wire __A08_NET_144;
    wire __A08_NET_145;
    wire __A08_NET_146;
    wire __A08_NET_147;
    wire __A08_NET_148;
    wire __A08_NET_150;
    wire __A08_NET_154;
    wire __A08_NET_155;
    wire __A08_NET_156;
    wire __A08_NET_157;
    wire __A08_NET_158;
    wire __A08_NET_159;
    wire __A08_NET_160;
    wire __A08_NET_161;
    wire __A08_NET_163;
    wire __A08_NET_164;
    wire __A08_NET_165;
    wire __A08_NET_171;
    wire __A08_NET_172;
    wire __A08_NET_173;
    wire __A08_NET_174;
    wire __A08_NET_175;
    wire __A08_NET_176;
    wire __A08_NET_177;
    wire __A08_NET_178;
    wire __A08_NET_179;
    wire __A08_NET_180;
    wire __A08_NET_181;
    wire __A08_NET_182;
    wire __A08_NET_183;
    wire __A08_NET_184;
    wire __A08_NET_185;
    wire __A08_NET_186;
    wire __A08_NET_187;
    wire __A08_NET_188;
    wire __A08_NET_189;
    wire __A08_NET_190;
    wire __A08_NET_191;
    wire __A08_NET_192;
    wire __A08_NET_193;
    wire __A08_NET_194;
    wire __A08_NET_195;
    wire __A08_NET_196;
    wire __A08_NET_197;
    wire __A08_NET_198;
    wire __A08_NET_203;
    wire __A08_NET_204;
    wire __A08_NET_205;
    wire __A08_NET_206;
    wire __A08_NET_207;
    wire __A08_NET_209;
    wire __A08_NET_210;
    wire __A08_NET_213;
    wire __A08_NET_214;
    wire __A08_NET_215;
    wire __A08_NET_216;
    wire __A08_NET_217;
    wire __A08_NET_218;
    wire __A08_NET_219;
    wire __A08_NET_220;
    wire __A08_NET_221;
    wire __A08_NET_222;
    wire __A08_NET_223;
    wire __A08_NET_224;
    wire __A08_NET_225;
    wire __A08_NET_226;
    wire __A08_NET_227;
    wire __A08_NET_228;
    wire __A08_NET_229;
    wire __A08_NET_230;
    wire __A08_NET_231;
    wire __A08_NET_232;
    wire __A08_NET_233;
    wire __A08_NET_234;
    wire __A08_NET_235;
    wire __A08_NET_236;
    wire __A08_NET_237;
    wire __A08_NET_238;
    wire __A08_NET_239;
    wire __A08_NET_240;
    wire __A08_NET_241;
    wire __A08_NET_243;
    wire __A08_NET_247;
    wire __A08_NET_248;
    wire __A08_NET_249;
    wire __A08_NET_250;
    wire __A08_NET_251;
    wire __A08_NET_252;
    wire __A08_NET_253;
    wire __A08_NET_254;
    wire __A08_NET_255;
    wire __A08_NET_257;
    wire __A08_NET_258;
    wire __A08_NET_265;
    wire __A08_NET_266;
    wire __A08_NET_267;
    wire __A08_NET_268;
    wire __A08_NET_269;
    wire __A08_NET_270;
    wire __A08_NET_271;
    wire __A08_NET_272;
    wire __A08_NET_273;
    wire __A08_NET_274;
    wire __A08_NET_275;
    wire __A08_NET_276;
    wire __A08_NET_277;
    wire __A08_NET_278;
    wire __A08_NET_279;
    wire __A08_NET_280;
    wire __A08_NET_281;
    wire __A08_NET_282;
    wire __A08_NET_283;
    wire __A08_NET_284;
    wire __A08_NET_285;
    wire __A08_NET_286;
    wire __A08_NET_287;
    wire __A08_NET_288;
    wire __A08_NET_289;
    wire __A08_NET_290;
    wire __A08_NET_291;
    wire __A08_NET_292;
    wire __A08_NET_293;
    wire __A08_NET_297;
    wire __A08_NET_298;
    wire __A08_NET_299;
    wire __A08_NET_300;
    wire __A08_NET_302;
    wire __A08_NET_303;
    wire __A08_NET_306;
    wire __A08_NET_307;
    wire __A08_NET_308;
    wire __A08_NET_309;
    wire __A08_NET_310;
    wire __A08_NET_311;
    wire __A08_NET_312;
    wire __A08_NET_313;
    wire __A08_NET_314;
    wire __A08_NET_315;
    wire __A08_NET_316;
    wire __A08_NET_317;
    wire __A08_NET_318;
    wire __A08_NET_319;
    wire __A08_NET_320;
    wire __A08_NET_321;
    wire __A08_NET_322;
    wire __A09_1__X1;
    wire __A09_1__X1_n;
    wire __A09_1__X2;
    wire __A09_1__X2_n;
    wire __A09_1__Y1;
    wire __A09_1__Y1_n;
    wire __A09_1__Y2;
    wire __A09_1__Y2_n;
    wire __A09_1___A1_n;
    wire __A09_1___A2_n;
    wire __A09_1___B1_n;
    wire __A09_1___B2_n;
    wire __A09_1___CI_INTERNAL;
    wire __A09_1___Q1_n;
    wire __A09_1___Q2_n;
    wire __A09_1___RL_OUT_1;
    wire __A09_1___RL_OUT_2;
    wire __A09_1___SUMA1;
    wire __A09_1___SUMA2;
    wire __A09_1___SUMB1;
    wire __A09_1___SUMB2;
    wire __A09_1___Z1_n;
    wire __A09_1___Z1_n_U9007_8;
    wire __A09_1___Z2_n;
    wire __A09_1___Z2_n_U9028_4;
    wire __A09_2__X1;
    wire __A09_2__X1_n;
    wire __A09_2__X2;
    wire __A09_2__X2_n;
    wire __A09_2__Y1;
    wire __A09_2__Y1_n;
    wire __A09_2__Y2;
    wire __A09_2__Y2_n;
    wire __A09_2___A1_n;
    wire __A09_2___A2_n;
    wire __A09_2___B1_n;
    wire __A09_2___B2_n;
    wire __A09_2___CI_INTERNAL;
    wire __A09_2___Q1_n;
    wire __A09_2___Q2_n;
    wire __A09_2___RL1_n;
    wire __A09_2___RL1_n_U9041_10;
    wire __A09_2___RL1_n_U9041_12;
    wire __A09_2___RL1_n_U9041_4;
    wire __A09_2___RL1_n_U9050_4;
    wire __A09_2___RL2_n;
    wire __A09_2___RL2_n_U9050_10;
    wire __A09_2___RL2_n_U9061_2;
    wire __A09_2___RL2_n_U9061_6;
    wire __A09_2___RL2_n_U9061_8;
    wire __A09_2___RL_OUT_1;
    wire __A09_2___RL_OUT_2;
    wire __A09_2___SUMA1;
    wire __A09_2___SUMA2;
    wire __A09_2___SUMB1;
    wire __A09_2___SUMB2;
    wire __A09_2___Z1_n;
    wire __A09_2___Z1_n_U9041_8;
    wire __A09_2___Z2_n;
    wire __A09_2___Z2_n_U9061_4;
    wire __A09_NET_130;
    wire __A09_NET_131;
    wire __A09_NET_132;
    wire __A09_NET_133;
    wire __A09_NET_134;
    wire __A09_NET_135;
    wire __A09_NET_136;
    wire __A09_NET_137;
    wire __A09_NET_138;
    wire __A09_NET_139;
    wire __A09_NET_140;
    wire __A09_NET_141;
    wire __A09_NET_143;
    wire __A09_NET_147;
    wire __A09_NET_148;
    wire __A09_NET_149;
    wire __A09_NET_150;
    wire __A09_NET_151;
    wire __A09_NET_152;
    wire __A09_NET_153;
    wire __A09_NET_154;
    wire __A09_NET_156;
    wire __A09_NET_157;
    wire __A09_NET_158;
    wire __A09_NET_164;
    wire __A09_NET_165;
    wire __A09_NET_166;
    wire __A09_NET_167;
    wire __A09_NET_168;
    wire __A09_NET_169;
    wire __A09_NET_170;
    wire __A09_NET_171;
    wire __A09_NET_172;
    wire __A09_NET_173;
    wire __A09_NET_174;
    wire __A09_NET_175;
    wire __A09_NET_176;
    wire __A09_NET_177;
    wire __A09_NET_178;
    wire __A09_NET_179;
    wire __A09_NET_180;
    wire __A09_NET_181;
    wire __A09_NET_182;
    wire __A09_NET_183;
    wire __A09_NET_184;
    wire __A09_NET_185;
    wire __A09_NET_186;
    wire __A09_NET_187;
    wire __A09_NET_188;
    wire __A09_NET_189;
    wire __A09_NET_190;
    wire __A09_NET_191;
    wire __A09_NET_196;
    wire __A09_NET_197;
    wire __A09_NET_198;
    wire __A09_NET_199;
    wire __A09_NET_200;
    wire __A09_NET_202;
    wire __A09_NET_203;
    wire __A09_NET_206;
    wire __A09_NET_207;
    wire __A09_NET_208;
    wire __A09_NET_209;
    wire __A09_NET_210;
    wire __A09_NET_211;
    wire __A09_NET_212;
    wire __A09_NET_213;
    wire __A09_NET_214;
    wire __A09_NET_215;
    wire __A09_NET_216;
    wire __A09_NET_217;
    wire __A09_NET_218;
    wire __A09_NET_219;
    wire __A09_NET_220;
    wire __A09_NET_221;
    wire __A09_NET_222;
    wire __A09_NET_223;
    wire __A09_NET_224;
    wire __A09_NET_225;
    wire __A09_NET_226;
    wire __A09_NET_227;
    wire __A09_NET_228;
    wire __A09_NET_229;
    wire __A09_NET_230;
    wire __A09_NET_231;
    wire __A09_NET_232;
    wire __A09_NET_233;
    wire __A09_NET_234;
    wire __A09_NET_236;
    wire __A09_NET_240;
    wire __A09_NET_241;
    wire __A09_NET_242;
    wire __A09_NET_243;
    wire __A09_NET_244;
    wire __A09_NET_245;
    wire __A09_NET_246;
    wire __A09_NET_247;
    wire __A09_NET_248;
    wire __A09_NET_250;
    wire __A09_NET_251;
    wire __A09_NET_258;
    wire __A09_NET_259;
    wire __A09_NET_260;
    wire __A09_NET_261;
    wire __A09_NET_262;
    wire __A09_NET_263;
    wire __A09_NET_264;
    wire __A09_NET_265;
    wire __A09_NET_266;
    wire __A09_NET_267;
    wire __A09_NET_268;
    wire __A09_NET_269;
    wire __A09_NET_270;
    wire __A09_NET_271;
    wire __A09_NET_272;
    wire __A09_NET_273;
    wire __A09_NET_274;
    wire __A09_NET_275;
    wire __A09_NET_276;
    wire __A09_NET_277;
    wire __A09_NET_278;
    wire __A09_NET_279;
    wire __A09_NET_280;
    wire __A09_NET_281;
    wire __A09_NET_282;
    wire __A09_NET_283;
    wire __A09_NET_284;
    wire __A09_NET_285;
    wire __A09_NET_286;
    wire __A09_NET_290;
    wire __A09_NET_291;
    wire __A09_NET_292;
    wire __A09_NET_293;
    wire __A09_NET_295;
    wire __A09_NET_296;
    wire __A09_NET_299;
    wire __A09_NET_300;
    wire __A09_NET_301;
    wire __A09_NET_302;
    wire __A09_NET_303;
    wire __A09_NET_304;
    wire __A09_NET_305;
    wire __A09_NET_306;
    wire __A09_NET_307;
    wire __A09_NET_308;
    wire __A09_NET_309;
    wire __A09_NET_310;
    wire __A09_NET_311;
    wire __A09_NET_312;
    wire __A09_NET_313;
    wire __A09_NET_314;
    wire __A09_NET_315;
    wire __A10_1__X1;
    wire __A10_1__X1_n;
    wire __A10_1__X2;
    wire __A10_1__X2_n;
    wire __A10_1__Y1;
    wire __A10_1__Y1_n;
    wire __A10_1__Y2;
    wire __A10_1__Y2_n;
    wire __A10_1___A1_n;
    wire __A10_1___A2_n;
    wire __A10_1___B1_n;
    wire __A10_1___B2_n;
    wire __A10_1___CI_INTERNAL;
    wire __A10_1___Q1_n;
    wire __A10_1___Q2_n;
    wire __A10_1___RL_OUT_1;
    wire __A10_1___RL_OUT_2;
    wire __A10_1___SUMA1;
    wire __A10_1___SUMA2;
    wire __A10_1___SUMB1;
    wire __A10_1___SUMB2;
    wire __A10_1___Z1_n;
    wire __A10_1___Z1_n_U10007_8;
    wire __A10_1___Z2_n;
    wire __A10_1___Z2_n_U10028_4;
    wire __A10_2__X1;
    wire __A10_2__X1_n;
    wire __A10_2__X2;
    wire __A10_2__X2_n;
    wire __A10_2__Y1;
    wire __A10_2__Y1_n;
    wire __A10_2__Y2;
    wire __A10_2__Y2_n;
    wire __A10_2___A1_n;
    wire __A10_2___A2_n;
    wire __A10_2___B1_n;
    wire __A10_2___B2_n;
    wire __A10_2___CI_INTERNAL;
    wire __A10_2___Q1_n;
    wire __A10_2___Q2_n;
    wire __A10_2___RL_OUT_1;
    wire __A10_2___RL_OUT_2;
    wire __A10_2___Z1_n;
    wire __A10_2___Z1_n_U10041_8;
    wire __A10_2___Z2_n;
    wire __A10_2___Z2_n_U10061_4;
    wire __A10_NET_129;
    wire __A10_NET_130;
    wire __A10_NET_131;
    wire __A10_NET_132;
    wire __A10_NET_133;
    wire __A10_NET_134;
    wire __A10_NET_135;
    wire __A10_NET_136;
    wire __A10_NET_137;
    wire __A10_NET_138;
    wire __A10_NET_139;
    wire __A10_NET_140;
    wire __A10_NET_142;
    wire __A10_NET_146;
    wire __A10_NET_147;
    wire __A10_NET_148;
    wire __A10_NET_149;
    wire __A10_NET_150;
    wire __A10_NET_151;
    wire __A10_NET_152;
    wire __A10_NET_153;
    wire __A10_NET_155;
    wire __A10_NET_156;
    wire __A10_NET_157;
    wire __A10_NET_163;
    wire __A10_NET_164;
    wire __A10_NET_165;
    wire __A10_NET_166;
    wire __A10_NET_167;
    wire __A10_NET_168;
    wire __A10_NET_169;
    wire __A10_NET_170;
    wire __A10_NET_171;
    wire __A10_NET_172;
    wire __A10_NET_173;
    wire __A10_NET_174;
    wire __A10_NET_175;
    wire __A10_NET_176;
    wire __A10_NET_177;
    wire __A10_NET_178;
    wire __A10_NET_179;
    wire __A10_NET_180;
    wire __A10_NET_181;
    wire __A10_NET_182;
    wire __A10_NET_183;
    wire __A10_NET_184;
    wire __A10_NET_185;
    wire __A10_NET_186;
    wire __A10_NET_187;
    wire __A10_NET_188;
    wire __A10_NET_189;
    wire __A10_NET_190;
    wire __A10_NET_195;
    wire __A10_NET_196;
    wire __A10_NET_197;
    wire __A10_NET_198;
    wire __A10_NET_199;
    wire __A10_NET_201;
    wire __A10_NET_202;
    wire __A10_NET_205;
    wire __A10_NET_206;
    wire __A10_NET_207;
    wire __A10_NET_208;
    wire __A10_NET_209;
    wire __A10_NET_210;
    wire __A10_NET_211;
    wire __A10_NET_212;
    wire __A10_NET_213;
    wire __A10_NET_214;
    wire __A10_NET_215;
    wire __A10_NET_216;
    wire __A10_NET_217;
    wire __A10_NET_218;
    wire __A10_NET_219;
    wire __A10_NET_220;
    wire __A10_NET_221;
    wire __A10_NET_222;
    wire __A10_NET_223;
    wire __A10_NET_224;
    wire __A10_NET_225;
    wire __A10_NET_226;
    wire __A10_NET_227;
    wire __A10_NET_228;
    wire __A10_NET_229;
    wire __A10_NET_230;
    wire __A10_NET_231;
    wire __A10_NET_232;
    wire __A10_NET_233;
    wire __A10_NET_235;
    wire __A10_NET_239;
    wire __A10_NET_240;
    wire __A10_NET_241;
    wire __A10_NET_242;
    wire __A10_NET_243;
    wire __A10_NET_244;
    wire __A10_NET_245;
    wire __A10_NET_246;
    wire __A10_NET_247;
    wire __A10_NET_249;
    wire __A10_NET_250;
    wire __A10_NET_257;
    wire __A10_NET_258;
    wire __A10_NET_259;
    wire __A10_NET_260;
    wire __A10_NET_261;
    wire __A10_NET_262;
    wire __A10_NET_263;
    wire __A10_NET_264;
    wire __A10_NET_265;
    wire __A10_NET_266;
    wire __A10_NET_267;
    wire __A10_NET_268;
    wire __A10_NET_269;
    wire __A10_NET_270;
    wire __A10_NET_271;
    wire __A10_NET_272;
    wire __A10_NET_273;
    wire __A10_NET_274;
    wire __A10_NET_275;
    wire __A10_NET_276;
    wire __A10_NET_277;
    wire __A10_NET_278;
    wire __A10_NET_279;
    wire __A10_NET_280;
    wire __A10_NET_281;
    wire __A10_NET_282;
    wire __A10_NET_283;
    wire __A10_NET_284;
    wire __A10_NET_285;
    wire __A10_NET_289;
    wire __A10_NET_290;
    wire __A10_NET_291;
    wire __A10_NET_292;
    wire __A10_NET_294;
    wire __A10_NET_295;
    wire __A10_NET_298;
    wire __A10_NET_299;
    wire __A10_NET_300;
    wire __A10_NET_301;
    wire __A10_NET_302;
    wire __A10_NET_303;
    wire __A10_NET_304;
    wire __A10_NET_305;
    wire __A10_NET_306;
    wire __A10_NET_307;
    wire __A10_NET_308;
    wire __A10_NET_309;
    wire __A10_NET_310;
    wire __A10_NET_311;
    wire __A10_NET_312;
    wire __A10_NET_313;
    wire __A10_NET_314;
    wire __A11_1__X1;
    wire __A11_1__X1_n;
    wire __A11_1__X2;
    wire __A11_1__X2_n;
    wire __A11_1__Y1;
    wire __A11_1__Y1_n;
    wire __A11_1__Y2;
    wire __A11_1__Y2_n;
    wire __A11_1___A1_n;
    wire __A11_1___A2_n;
    wire __A11_1___B1_n;
    wire __A11_1___B2_n;
    wire __A11_1___CI_INTERNAL;
    wire __A11_1___Q1_n;
    wire __A11_1___Q2_n;
    wire __A11_1___RL_OUT_1;
    wire __A11_1___RL_OUT_2;
    wire __A11_1___Z1_n;
    wire __A11_1___Z1_n_U11007_8;
    wire __A11_1___Z2_n;
    wire __A11_1___Z2_n_U11028_4;
    wire __A11_2__X1;
    wire __A11_2__X1_n;
    wire __A11_2__X2;
    wire __A11_2__X2_n;
    wire __A11_2__Y1;
    wire __A11_2__Y1_n;
    wire __A11_2__Y2;
    wire __A11_2__Y2_n;
    wire __A11_2___B1_n;
    wire __A11_2___B2_n;
    wire __A11_2___CI_INTERNAL;
    wire __A11_2___CO_OUT;
    wire __A11_2___CO_OUT_U11041_2;
    wire __A11_2___CO_OUT_U11050_2;
    wire __A11_2___GEM1;
    wire __A11_2___Q1_n;
    wire __A11_2___Q2_n;
    wire __A11_2___RL_OUT_1;
    wire __A11_NET_130;
    wire __A11_NET_131;
    wire __A11_NET_132;
    wire __A11_NET_133;
    wire __A11_NET_134;
    wire __A11_NET_135;
    wire __A11_NET_136;
    wire __A11_NET_137;
    wire __A11_NET_138;
    wire __A11_NET_139;
    wire __A11_NET_140;
    wire __A11_NET_141;
    wire __A11_NET_143;
    wire __A11_NET_147;
    wire __A11_NET_148;
    wire __A11_NET_149;
    wire __A11_NET_150;
    wire __A11_NET_151;
    wire __A11_NET_152;
    wire __A11_NET_153;
    wire __A11_NET_154;
    wire __A11_NET_156;
    wire __A11_NET_157;
    wire __A11_NET_158;
    wire __A11_NET_164;
    wire __A11_NET_165;
    wire __A11_NET_166;
    wire __A11_NET_167;
    wire __A11_NET_168;
    wire __A11_NET_169;
    wire __A11_NET_170;
    wire __A11_NET_171;
    wire __A11_NET_172;
    wire __A11_NET_173;
    wire __A11_NET_174;
    wire __A11_NET_175;
    wire __A11_NET_176;
    wire __A11_NET_177;
    wire __A11_NET_178;
    wire __A11_NET_179;
    wire __A11_NET_180;
    wire __A11_NET_181;
    wire __A11_NET_182;
    wire __A11_NET_183;
    wire __A11_NET_184;
    wire __A11_NET_185;
    wire __A11_NET_186;
    wire __A11_NET_187;
    wire __A11_NET_188;
    wire __A11_NET_189;
    wire __A11_NET_190;
    wire __A11_NET_191;
    wire __A11_NET_196;
    wire __A11_NET_197;
    wire __A11_NET_198;
    wire __A11_NET_199;
    wire __A11_NET_200;
    wire __A11_NET_202;
    wire __A11_NET_203;
    wire __A11_NET_206;
    wire __A11_NET_207;
    wire __A11_NET_208;
    wire __A11_NET_209;
    wire __A11_NET_210;
    wire __A11_NET_211;
    wire __A11_NET_212;
    wire __A11_NET_213;
    wire __A11_NET_214;
    wire __A11_NET_215;
    wire __A11_NET_216;
    wire __A11_NET_217;
    wire __A11_NET_218;
    wire __A11_NET_219;
    wire __A11_NET_220;
    wire __A11_NET_221;
    wire __A11_NET_222;
    wire __A11_NET_223;
    wire __A11_NET_224;
    wire __A11_NET_225;
    wire __A11_NET_226;
    wire __A11_NET_227;
    wire __A11_NET_228;
    wire __A11_NET_229;
    wire __A11_NET_230;
    wire __A11_NET_231;
    wire __A11_NET_232;
    wire __A11_NET_233;
    wire __A11_NET_234;
    wire __A11_NET_236;
    wire __A11_NET_240;
    wire __A11_NET_241;
    wire __A11_NET_242;
    wire __A11_NET_243;
    wire __A11_NET_244;
    wire __A11_NET_245;
    wire __A11_NET_246;
    wire __A11_NET_247;
    wire __A11_NET_248;
    wire __A11_NET_250;
    wire __A11_NET_251;
    wire __A11_NET_258;
    wire __A11_NET_259;
    wire __A11_NET_260;
    wire __A11_NET_261;
    wire __A11_NET_262;
    wire __A11_NET_263;
    wire __A11_NET_264;
    wire __A11_NET_265;
    wire __A11_NET_266;
    wire __A11_NET_267;
    wire __A11_NET_268;
    wire __A11_NET_269;
    wire __A11_NET_270;
    wire __A11_NET_271;
    wire __A11_NET_272;
    wire __A11_NET_273;
    wire __A11_NET_274;
    wire __A11_NET_275;
    wire __A11_NET_276;
    wire __A11_NET_277;
    wire __A11_NET_278;
    wire __A11_NET_279;
    wire __A11_NET_280;
    wire __A11_NET_281;
    wire __A11_NET_282;
    wire __A11_NET_283;
    wire __A11_NET_284;
    wire __A11_NET_285;
    wire __A11_NET_286;
    wire __A11_NET_290;
    wire __A11_NET_291;
    wire __A11_NET_292;
    wire __A11_NET_293;
    wire __A11_NET_295;
    wire __A11_NET_296;
    wire __A11_NET_299;
    wire __A11_NET_300;
    wire __A11_NET_301;
    wire __A11_NET_302;
    wire __A11_NET_303;
    wire __A11_NET_304;
    wire __A11_NET_305;
    wire __A11_NET_306;
    wire __A11_NET_307;
    wire __A11_NET_308;
    wire __A11_NET_309;
    wire __A11_NET_310;
    wire __A11_NET_311;
    wire __A11_NET_312;
    wire __A11_NET_313;
    wire __A11_NET_314;
    wire __A11_NET_315;
    wire __A12_1__G01A_n;
    wire __A12_1__G02_n;
    wire __A12_1__G03_n;
    wire __A12_1__G16A_n;
    wire __A12_1__GNZRO;
    wire __A12_1__GNZRO_U12016_2;
    wire __A12_1__GNZRO_U12016_4;
    wire __A12_1__PA03;
    wire __A12_1__PA03_n;
    wire __A12_1__PA06;
    wire __A12_1__PA06_n;
    wire __A12_1__PA09;
    wire __A12_1__PA09_n;
    wire __A12_1__PA12;
    wire __A12_1__PA12_n;
    wire __A12_1__PA15;
    wire __A12_1__PA15_n;
    wire __A12_1__PB09;
    wire __A12_1__PB09_n;
    wire __A12_1__PB15;
    wire __A12_1__PB15_n;
    wire __A12_1__PC15;
    wire __A12_1__T7PHS4;
    wire __A12_1__T7PHS4_n;
    wire __A12_2__G01A;
    wire __A12_NET_112;
    wire __A12_NET_113;
    wire __A12_NET_114;
    wire __A12_NET_115;
    wire __A12_NET_117;
    wire __A12_NET_118;
    wire __A12_NET_119;
    wire __A12_NET_120;
    wire __A12_NET_121;
    wire __A12_NET_122;
    wire __A12_NET_123;
    wire __A12_NET_124;
    wire __A12_NET_125;
    wire __A12_NET_126;
    wire __A12_NET_127;
    wire __A12_NET_128;
    wire __A12_NET_129;
    wire __A12_NET_130;
    wire __A12_NET_131;
    wire __A12_NET_132;
    wire __A12_NET_133;
    wire __A12_NET_134;
    wire __A12_NET_135;
    wire __A12_NET_136;
    wire __A12_NET_137;
    wire __A12_NET_138;
    wire __A12_NET_139;
    wire __A12_NET_140;
    wire __A12_NET_141;
    wire __A12_NET_142;
    wire __A12_NET_143;
    wire __A12_NET_149;
    wire __A12_NET_151;
    wire __A12_NET_153;
    wire __A12_NET_160;
    wire __A12_NET_161;
    wire __A12_NET_162;
    wire __A12_NET_167;
    wire __A12_NET_168;
    wire __A12_NET_171;
    wire __A12_NET_173;
    wire __A12_NET_178;
    wire __A12_NET_179;
    wire __A12_NET_180;
    wire __A12_NET_183;
    wire __A12_NET_184;
    wire __A12_NET_185;
    wire __A12_NET_187;
    wire __A12_NET_188;
    wire __A12_NET_189;
    wire __A12_NET_190;
    wire __A12_NET_191;
    wire __A12_NET_192;
    wire __A12_NET_195;
    wire __A12_NET_198;
    wire __A12_NET_199;
    wire __A12_NET_200;
    wire __A12_NET_201;
    wire __A12_NET_202;
    wire __A12_NET_203;
    wire __A12_NET_204;
    wire __A12_NET_205;
    wire __A12_NET_206;
    wire __A12_NET_207;
    wire __A12_NET_208;
    wire __A12_NET_209;
    wire __A12_NET_210;
    wire __A12_NET_211;
    wire __A12_NET_212;
    wire __A12_NET_213;
    wire __A12_NET_214;
    wire __A12_NET_215;
    wire __A12_NET_216;
    wire __A12_NET_217;
    wire __A12_NET_218;
    wire __A12_NET_219;
    wire __A12_NET_220;
    wire __A12_NET_221;
    wire __A12_NET_222;
    wire __A12_NET_223;
    wire __A12_NET_225;
    wire __A12_NET_226;
    wire __A12_NET_227;
    wire __A12_NET_228;
    wire __A12_NET_229;
    wire __A12_NET_230;
    wire __A12_NET_231;
    wire __A12_NET_232;
    wire __A12_NET_233;
    wire __A12_NET_234;
    wire __A12_NET_236;
    wire __A12_NET_237;
    wire __A12_NET_238;
    wire __A12_NET_239;
    wire __A12_NET_240;
    wire __A12_NET_241;
    wire __A12_NET_243;
    wire __A12_NET_244;
    wire __A12_NET_245;
    wire __A12_NET_246;
    wire __A12_NET_247;
    wire __A12_NET_248;
    wire __A12_NET_249;
    wire __A12_NET_250;
    wire __A12_NET_251;
    wire __A12_NET_252;
    wire __A12_NET_253;
    wire __A12_NET_254;
    wire __A12_NET_255;
    wire __A12_NET_256;
    wire __A12_NET_257;
    wire __A13_1__CGCWAR;
    wire __A13_1__CKTAL_n;
    wire __A13_1__CKTAL_n_U13006_2;
    wire __A13_1__CKTAL_n_U13006_4;
    wire __A13_1__CON1;
    wire __A13_1__CON2;
    wire __A13_1__CON3;
    wire __A13_1__DOFILT;
    wire __A13_1__F12B_n;
    wire __A13_1__F14H;
    wire __A13_1__FILTIN;
    wire __A13_1__FS13_n;
    wire __A13_1__NOTEST;
    wire __A13_1__NOTEST_n;
    wire __A13_1__SBYEXT;
    wire __A13_1__SCADBL;
    wire __A13_1__SCAS10;
    wire __A13_1__SCAS17;
    wire __A13_1__SYNC14_n;
    wire __A13_1__SYNC4_n;
    wire __A13_1__TEMPIN_n;
    wire __A13_1__WARN;
    wire __A13_1__WATCH;
    wire __A13_1__WATCHP;
    wire __A13_2__INOTRD;
    wire __A13_2__STORE1;
    wire __A13_NET_164;
    wire __A13_NET_165;
    wire __A13_NET_166;
    wire __A13_NET_167;
    wire __A13_NET_170;
    wire __A13_NET_171;
    wire __A13_NET_172;
    wire __A13_NET_174;
    wire __A13_NET_175;
    wire __A13_NET_176;
    wire __A13_NET_177;
    wire __A13_NET_178;
    wire __A13_NET_179;
    wire __A13_NET_179_U13121_2;
    wire __A13_NET_179_U13121_4;
    wire __A13_NET_180;
    wire __A13_NET_183;
    wire __A13_NET_184;
    wire __A13_NET_186;
    wire __A13_NET_187;
    wire __A13_NET_188;
    wire __A13_NET_189;
    wire __A13_NET_190;
    wire __A13_NET_191;
    wire __A13_NET_192;
    wire __A13_NET_195;
    wire __A13_NET_196;
    wire __A13_NET_197;
    wire __A13_NET_198;
    wire __A13_NET_201;
    wire __A13_NET_204;
    wire __A13_NET_205;
    wire __A13_NET_206;
    wire __A13_NET_207;
    wire __A13_NET_211;
    wire __A13_NET_212;
    wire __A13_NET_213;
    wire __A13_NET_215;
    wire __A13_NET_216;
    wire __A13_NET_217;
    wire __A13_NET_220;
    wire __A13_NET_221;
    wire __A13_NET_227;
    wire __A13_NET_228;
    wire __A13_NET_231;
    wire __A13_NET_232;
    wire __A13_NET_233;
    wire __A13_NET_234;
    wire __A13_NET_235;
    wire __A13_NET_236;
    wire __A13_NET_237;
    wire __A13_NET_238;
    wire __A13_NET_241;
    wire __A13_NET_242;
    wire __A13_NET_243;
    wire __A13_NET_248;
    wire __A13_NET_251;
    wire __A13_NET_252;
    wire __A13_NET_253;
    wire __A13_NET_254;
    wire __A13_NET_255;
    wire __A13_NET_256;
    wire __A13_NET_257;
    wire __A13_NET_260;
    wire __A13_NET_261;
    wire __A13_NET_262;
    wire __A13_NET_264;
    wire __A13_NET_266;
    wire __A13_NET_267;
    wire __A13_NET_268;
    wire __A13_NET_270;
    wire __A13_NET_271;
    wire __A13_NET_272;
    wire __A13_NET_273;
    wire __A13_NET_274;
    wire __A13_NET_277;
    wire __A13_NET_277_U13006_10;
    wire __A13_NET_277_U13006_12;
    wire __A13_NET_277_U13006_6;
    wire __A13_NET_277_U13006_8;
    wire __A13_NET_277_U13036_12;
    wire __A13_NET_277_U13036_2;
    wire __A13_NET_277_U13036_4;
    wire __A13_NET_277_U13036_6;
    wire __A13_NET_277_U13051_2;
    wire __A13_NET_277_U13051_4;
    wire __A13_NET_277_U13051_6;
    wire __A13_NET_278;
    wire __A13_NET_279;
    wire __A13_NET_280;
    wire __A13_NET_281;
    wire __A13_NET_282;
    wire __A13_NET_283;
    wire __A13_NET_284;
    wire __A13_NET_285;
    wire __A13_NET_286;
    wire __A13_NET_287;
    wire __A13_NET_290;
    wire __A13_NET_291;
    wire __A13_NET_292;
    wire __A13_NET_293;
    wire __A13_NET_294;
    wire __A13_NET_295;
    wire __A13_NET_297;
    wire __A13_NET_301;
    wire __A13_NET_302;
    wire __A13_NET_303;
    wire __A13_NET_304;
    wire __A13_NET_305;
    wire __A13_NET_306;
    wire __A13_NET_307;
    wire __A13_NET_307_U13036_10;
    wire __A13_NET_307_U13036_8;
    wire __A13_NET_308;
    wire __A13_NET_309;
    wire __A13_NET_310;
    wire __A13_NET_311;
    wire __A13_NET_312;
    wire __A13_NET_313;
    wire __A13_NET_314;
    wire __A13_NET_315;
    wire __A13_NET_316;
    wire __A13_NET_317;
    wire __A13_NET_318;
    wire __A13_NET_319;
    wire __A13_NET_320;
    wire __A13_NET_321;
    wire __A13_NET_322;
    wire __A13_NET_323;
    wire __A13_NET_324;
    wire __A14_1__CLEARA;
    wire __A14_1__CLEARB;
    wire __A14_1__CLEARC;
    wire __A14_1__CLEARD;
    wire __A14_1__ERAS;
    wire __A14_1__ERAS_U14014_10;
    wire __A14_1__ERAS_U14014_12;
    wire __A14_1__ERAS_n;
    wire __A14_1__FNERAS_n;
    wire __A14_1__IHENV;
    wire __A14_1__REDRST;
    wire __A14_1__ROP_n;
    wire __A14_1__RSTK_n;
    wire __A14_1__S08A;
    wire __A14_1__S08A_n;
    wire __A14_1__SBESET;
    wire __A14_1__SBFSET;
    wire __A14_1__SBFSET_U14014_2;
    wire __A14_1__SBFSET_U14014_4;
    wire __A14_1__SETAB_n;
    wire __A14_1__SETCD_n;
    wire __A14_1__TPGE;
    wire __A14_1__TPGE_U14033_2;
    wire __A14_1__TPGE_U14033_4;
    wire __A14_1__TPGF;
    wire __A14_1__TPGF_U14014_6;
    wire __A14_1__TPGF_U14014_8;
    wire __A14_2__EAD09;
    wire __A14_2__EAD09_n;
    wire __A14_2__EAD10;
    wire __A14_2__EAD10_n;
    wire __A14_2__EAD11;
    wire __A14_2__EAD11_n;
    wire __A14_2__IL01_n;
    wire __A14_2__IL02_n;
    wire __A14_2__IL03_n;
    wire __A14_2__IL04_n;
    wire __A14_2__IL05_n;
    wire __A14_2__IL06_n;
    wire __A14_2__IL07_n;
    wire __A14_2__ILP;
    wire __A14_2__ILP_n;
    wire __A14_2__RILP1;
    wire __A14_2__RILP1_n;
    wire __A14_2__XB0E;
    wire __A14_2__XT0;
    wire __A14_2__XT0E;
    wire __A14_2__XT1;
    wire __A14_2__XT2;
    wire __A14_2__XT3;
    wire __A14_2__XT4;
    wire __A14_2__XT5;
    wire __A14_2__XT6;
    wire __A14_2__XT7;
    wire __A14_2__XT7_n;
    wire __A14_2__YB0;
    wire __A14_2__YB0E;
    wire __A14_2__YB1;
    wire __A14_2__YB1_n;
    wire __A14_2__YB2;
    wire __A14_2__YB2_n;
    wire __A14_2__YB3;
    wire __A14_2__YB3_n;
    wire __A14_2__YT0;
    wire __A14_2__YT0E;
    wire __A14_2__YT1;
    wire __A14_2__YT1_n;
    wire __A14_2__YT2;
    wire __A14_2__YT2_n;
    wire __A14_2__YT3;
    wire __A14_2__YT3_n;
    wire __A14_2__YT4;
    wire __A14_2__YT4_n;
    wire __A14_2__YT5;
    wire __A14_2__YT5_n;
    wire __A14_2__YT6;
    wire __A14_2__YT6_n;
    wire __A14_2__YT7;
    wire __A14_2__YT7_n;
    wire __A14_NET_192;
    wire __A14_NET_193;
    wire __A14_NET_194;
    wire __A14_NET_195;
    wire __A14_NET_196;
    wire __A14_NET_197;
    wire __A14_NET_198;
    wire __A14_NET_199;
    wire __A14_NET_200;
    wire __A14_NET_201;
    wire __A14_NET_202;
    wire __A14_NET_203;
    wire __A14_NET_204;
    wire __A14_NET_205;
    wire __A14_NET_206;
    wire __A14_NET_207;
    wire __A14_NET_208;
    wire __A14_NET_209;
    wire __A14_NET_210;
    wire __A14_NET_211;
    wire __A14_NET_212;
    wire __A14_NET_213;
    wire __A14_NET_214;
    wire __A14_NET_215;
    wire __A14_NET_216;
    wire __A14_NET_217;
    wire __A14_NET_219;
    wire __A14_NET_220;
    wire __A14_NET_221;
    wire __A14_NET_223;
    wire __A14_NET_224;
    wire __A14_NET_227;
    wire __A14_NET_228;
    wire __A14_NET_229;
    wire __A14_NET_230;
    wire __A14_NET_231;
    wire __A14_NET_232;
    wire __A14_NET_233;
    wire __A14_NET_234;
    wire __A14_NET_235;
    wire __A14_NET_236;
    wire __A14_NET_237;
    wire __A14_NET_238;
    wire __A14_NET_239;
    wire __A14_NET_240;
    wire __A14_NET_241;
    wire __A14_NET_242;
    wire __A14_NET_243;
    wire __A14_NET_244;
    wire __A14_NET_245;
    wire __A14_NET_248;
    wire __A14_NET_249;
    wire __A14_NET_251;
    wire __A14_NET_252;
    wire __A14_NET_253;
    wire __A14_NET_254;
    wire __A14_NET_256;
    wire __A14_NET_257;
    wire __A14_NET_258;
    wire __A14_NET_259;
    wire __A14_NET_260;
    wire __A14_NET_261;
    wire __A14_NET_262;
    wire __A14_NET_263;
    wire __A14_NET_264;
    wire __A14_NET_265;
    wire __A14_NET_266;
    wire __A14_NET_267;
    wire __A14_NET_268;
    wire __A14_NET_269;
    wire __A14_NET_270;
    wire __A14_NET_273;
    wire __A14_NET_274;
    wire __A14_NET_279;
    wire __A14_NET_280;
    wire __A14_NET_285;
    wire __A14_NET_286;
    wire __A14_NET_290;
    wire __A14_NET_291;
    wire __A14_NET_292;
    wire __A14_NET_294;
    wire __A14_NET_295;
    wire __A14_NET_296;
    wire __A14_NET_298;
    wire __A14_NET_299;
    wire __A14_NET_300;
    wire __A14_NET_301;
    wire __A14_NET_302;
    wire __A14_NET_305;
    wire __A15_1__BBK1;
    wire __A15_1__BBK2;
    wire __A15_1__BBK3;
    wire __A15_1__BK16;
    wire __A15_1__DNRPTA;
    wire __A15_1__EB10_n;
    wire __A15_1__EB11;
    wire __A15_1__EB9_n;
    wire __A15_1__F11;
    wire __A15_1__F11_n;
    wire __A15_1__F12;
    wire __A15_1__F12_n;
    wire __A15_1__F13;
    wire __A15_1__F13_n;
    wire __A15_1__F14;
    wire __A15_1__F14_n;
    wire __A15_1__F15;
    wire __A15_1__F15_n;
    wire __A15_1__F16;
    wire __A15_1__F16_n;
    wire __A15_1__FB11;
    wire __A15_1__FB11_n;
    wire __A15_1__FB12;
    wire __A15_1__FB12_n;
    wire __A15_1__FB13;
    wire __A15_1__FB13_n;
    wire __A15_1__FB14;
    wire __A15_1__FB14_n;
    wire __A15_1__FB16;
    wire __A15_1__FB16_n;
    wire __A15_1__KRPTA_n;
    wire __A15_1__PRPOR1;
    wire __A15_1__PRPOR2;
    wire __A15_1__PRPOR3;
    wire __A15_1__PRPOR4;
    wire __A15_1__RPTA12;
    wire __A15_1__RPTAD6;
    wire __A15_1__RRPA1_n;
    wire __A15_2__036H;
    wire __A15_2__036L;
    wire __A15_2__147H;
    wire __A15_2__147L;
    wire __A15_2__2510H;
    wire __A15_2__2510L;
    wire __A15_2__KY1RST;
    wire __A15_2__KY2RST;
    wire __A15_2__NE00;
    wire __A15_2__NE01;
    wire __A15_2__NE012_n;
    wire __A15_2__NE02;
    wire __A15_2__NE03;
    wire __A15_2__NE036_n;
    wire __A15_2__NE04;
    wire __A15_2__NE05;
    wire __A15_2__NE06;
    wire __A15_2__NE07;
    wire __A15_2__NE10;
    wire __A15_2__NE147_n;
    wire __A15_2__NE2510_n;
    wire __A15_2__NE345_n;
    wire __A15_2__NE6710_n;
    wire __A15_2__RPTAD3;
    wire __A15_2__RPTAD4;
    wire __A15_2__RPTAD5;
    wire __A15_NET_149;
    wire __A15_NET_150;
    wire __A15_NET_151;
    wire __A15_NET_152;
    wire __A15_NET_153;
    wire __A15_NET_154;
    wire __A15_NET_155;
    wire __A15_NET_156;
    wire __A15_NET_157;
    wire __A15_NET_158;
    wire __A15_NET_159;
    wire __A15_NET_160;
    wire __A15_NET_161;
    wire __A15_NET_162;
    wire __A15_NET_163;
    wire __A15_NET_164;
    wire __A15_NET_165;
    wire __A15_NET_166;
    wire __A15_NET_167;
    wire __A15_NET_168;
    wire __A15_NET_171;
    wire __A15_NET_174;
    wire __A15_NET_175;
    wire __A15_NET_176;
    wire __A15_NET_177;
    wire __A15_NET_179;
    wire __A15_NET_181;
    wire __A15_NET_184;
    wire __A15_NET_185;
    wire __A15_NET_186;
    wire __A15_NET_187;
    wire __A15_NET_188;
    wire __A15_NET_189;
    wire __A15_NET_192;
    wire __A15_NET_195;
    wire __A15_NET_197;
    wire __A15_NET_198;
    wire __A15_NET_199;
    wire __A15_NET_200;
    wire __A15_NET_201;
    wire __A15_NET_202;
    wire __A15_NET_203;
    wire __A15_NET_204;
    wire __A15_NET_205;
    wire __A15_NET_206;
    wire __A15_NET_207;
    wire __A15_NET_208;
    wire __A15_NET_209;
    wire __A15_NET_210;
    wire __A15_NET_213;
    wire __A15_NET_214;
    wire __A15_NET_215;
    wire __A15_NET_216;
    wire __A15_NET_217;
    wire __A15_NET_218;
    wire __A15_NET_219;
    wire __A15_NET_220;
    wire __A15_NET_221;
    wire __A15_NET_222;
    wire __A15_NET_223;
    wire __A15_NET_224;
    wire __A15_NET_225;
    wire __A15_NET_226;
    wire __A15_NET_227;
    wire __A15_NET_228;
    wire __A15_NET_229;
    wire __A15_NET_229_U15016_10;
    wire __A15_NET_229_U15016_8;
    wire __A15_NET_232;
    wire __A15_NET_232_U15016_12;
    wire __A15_NET_232_U15039_2;
    wire __A15_NET_234;
    wire __A15_NET_235;
    wire __A15_NET_236;
    wire __A15_NET_237;
    wire __A15_NET_238;
    wire __A15_NET_239;
    wire __A15_NET_240;
    wire __A15_NET_241;
    wire __A15_NET_242;
    wire __A15_NET_243;
    wire __A15_NET_244;
    wire __A15_NET_245;
    wire __A15_NET_246;
    wire __A15_NET_251;
    wire __A15_NET_260;
    wire __A15_NET_261;
    wire __A15_NET_262;
    wire __A15_NET_265;
    wire __A15_NET_266;
    wire __A15_NET_267;
    wire __A15_NET_268;
    wire __A15_NET_269;
    wire __A15_NET_270;
    wire __A15_NET_271;
    wire __A15_NET_272;
    wire __A15_NET_273;
    wire __A15_NET_274;
    wire __A15_NET_282;
    wire __A15_NET_283;
    wire __A15_NET_284;
    wire __A15_NET_285;
    wire __A15_NET_286;
    wire __A15_NET_287;
    wire __A15_NET_290;
    wire __A15_NET_291;
    wire __A15_NET_294;
    wire __A15_NET_295;
    wire __A15_NET_296;
    wire __A15_NET_297;
    wire __A15_NET_298;
    wire __A15_NET_299;
    wire __A15_NET_300;
    wire __A15_NET_301;
    wire __A15_NET_302;
    wire __A15_NET_303;
    wire __A15_NET_304;
    wire __A15_NET_305;
    wire __A15_NET_306;
    wire __A15_NET_307;
    wire __A15_NET_310;
    wire __A16_1__CCH05;
    wire __A16_1__CCH06;
    wire __A16_1__CH1207;
    wire __A16_1__OT1207;
    wire __A16_1__OT1207_n;
    wire __A16_1__RCH05_n;
    wire __A16_1__RCH06_n;
    wire __A16_1__RCmXmP;
    wire __A16_1__RCmXmY;
    wire __A16_1__RCmXpP;
    wire __A16_1__RCmXpY;
    wire __A16_1__RCmYmR;
    wire __A16_1__RCmYpR;
    wire __A16_1__RCmZmR;
    wire __A16_1__RCmZpR;
    wire __A16_1__RCpXmP;
    wire __A16_1__RCpXmY;
    wire __A16_1__RCpXpP;
    wire __A16_1__RCpXpY;
    wire __A16_1__RCpYmR;
    wire __A16_1__RCpYpR;
    wire __A16_1__RCpZmR;
    wire __A16_1__RCpZpR;
    wire __A16_1__TVCNAB;
    wire __A16_1__WCH05_n;
    wire __A16_1__WCH06_n;
    wire __A16_2__COARSE;
    wire __A16_2__DISDAC;
    wire __A16_2__ENERIM;
    wire __A16_2__ENEROP;
    wire __A16_2__ISSWAR;
    wire __A16_2__MROLGT;
    wire __A16_2__S4BOFF;
    wire __A16_2__S4BSEQ;
    wire __A16_2__S4BTAK;
    wire __A16_2__STARON;
    wire __A16_2__ZEROPT;
    wire __A16_2__ZIMCDU;
    wire __A16_2__ZOPCDU;
    wire __A16_NET_102;
    wire __A16_NET_103;
    wire __A16_NET_104;
    wire __A16_NET_105;
    wire __A16_NET_106;
    wire __A16_NET_107;
    wire __A16_NET_108;
    wire __A16_NET_109;
    wire __A16_NET_110;
    wire __A16_NET_111;
    wire __A16_NET_112;
    wire __A16_NET_113;
    wire __A16_NET_114;
    wire __A16_NET_115;
    wire __A16_NET_116;
    wire __A16_NET_117;
    wire __A16_NET_118;
    wire __A16_NET_119;
    wire __A16_NET_120;
    wire __A16_NET_121;
    wire __A16_NET_122;
    wire __A16_NET_123;
    wire __A16_NET_124;
    wire __A16_NET_125;
    wire __A16_NET_126;
    wire __A16_NET_127;
    wire __A16_NET_128;
    wire __A16_NET_129;
    wire __A16_NET_130;
    wire __A16_NET_131;
    wire __A16_NET_132;
    wire __A16_NET_133;
    wire __A16_NET_134;
    wire __A16_NET_135;
    wire __A16_NET_136;
    wire __A16_NET_137;
    wire __A16_NET_138;
    wire __A16_NET_139;
    wire __A16_NET_140;
    wire __A16_NET_141;
    wire __A16_NET_142;
    wire __A16_NET_143;
    wire __A16_NET_144;
    wire __A16_NET_145;
    wire __A16_NET_146;
    wire __A16_NET_147;
    wire __A16_NET_148;
    wire __A16_NET_149;
    wire __A16_NET_150;
    wire __A16_NET_151;
    wire __A16_NET_152;
    wire __A16_NET_153;
    wire __A16_NET_154;
    wire __A16_NET_155;
    wire __A16_NET_156;
    wire __A16_NET_157;
    wire __A16_NET_159;
    wire __A16_NET_160;
    wire __A16_NET_163;
    wire __A16_NET_164;
    wire __A16_NET_165;
    wire __A16_NET_166;
    wire __A16_NET_167;
    wire __A16_NET_168;
    wire __A16_NET_169;
    wire __A16_NET_170;
    wire __A16_NET_171;
    wire __A16_NET_172;
    wire __A16_NET_173;
    wire __A16_NET_174;
    wire __A16_NET_175;
    wire __A16_NET_176;
    wire __A16_NET_177;
    wire __A16_NET_178;
    wire __A16_NET_179;
    wire __A16_NET_180;
    wire __A16_NET_181;
    wire __A16_NET_182;
    wire __A16_NET_183;
    wire __A16_NET_184;
    wire __A16_NET_185;
    wire __A16_NET_186;
    wire __A16_NET_187;
    wire __A16_NET_191;
    wire __A16_NET_192;
    wire __A16_NET_193;
    wire __A16_NET_194;
    wire __A16_NET_195;
    wire __A16_NET_196;
    wire __A16_NET_197;
    wire __A16_NET_198;
    wire __A16_NET_199;
    wire __A16_NET_200;
    wire __A16_NET_201;
    wire __A16_NET_202;
    wire __A16_NET_203;
    wire __A16_NET_204;
    wire __A16_NET_205;
    wire __A16_NET_206;
    wire __A16_NET_207;
    wire __A16_NET_208;
    wire __A16_NET_209;
    wire __A16_NET_210;
    wire __A16_NET_211;
    wire __A16_NET_212;
    wire __A16_NET_213;
    wire __A16_NET_214;
    wire __A16_NET_215;
    wire __A16_NET_216;
    wire __A16_NET_217;
    wire __A16_NET_218;
    wire __A16_NET_219;
    wire __A16_NET_220;
    wire __A16_NET_221;
    wire __A16_NET_222;
    wire __A16_NET_223;
    wire __A16_NET_224;
    wire __A16_NET_225;
    wire __A16_NET_226;
    wire __A16_NET_227;
    wire __A16_NET_228;
    wire __A16_NET_229;
    wire __A16_NET_230;
    wire __A16_NET_231;
    wire __A16_NET_232;
    wire __A16_NET_233;
    wire __A16_NET_234;
    wire __A16_NET_235;
    wire __A16_NET_236;
    wire __A16_NET_237;
    wire __A16_NET_238;
    wire __A16_NET_239;
    wire __A16_NET_240;
    wire __A16_NET_241;
    wire __A16_NET_242;
    wire __A16_NET_243;
    wire __A16_NET_244;
    wire __A16_NET_245;
    wire __A16_NET_246;
    wire __A16_NET_247;
    wire __A16_NET_248;
    wire __A16_NET_249;
    wire __A16_NET_250;
    wire __A16_NET_251;
    wire __A16_NET_252;
    wire __A16_NET_253;
    wire __A16_NET_254;
    wire __A16_NET_255;
    wire __A16_NET_256;
    wire __A16_NET_257;
    wire __A16_NET_258;
    wire __A16_NET_259;
    wire __A16_NET_260;
    wire __A16_NET_261;
    wire __A16_NET_262;
    wire __A16_NET_263;
    wire __A16_NET_264;
    wire __A16_NET_265;
    wire __A16_NET_266;
    wire __A16_NET_267;
    wire __A16_NET_268;
    wire __A16_NET_269;
    wire __A16_NET_270;
    wire __A16_NET_271;
    wire __A16_NET_272;
    wire __A16_NET_273;
    wire __A16_NET_274;
    wire __A17_1__F04B_n;
    wire __A17_1__FO5D;
    wire __A17_1__RCH30_n;
    wire __A17_1__RCH31_n;
    wire __A17_1__RCH32_n;
    wire __A17_1__TRP31A;
    wire __A17_1__TRP31B;
    wire __A17_1__TRP32;
    wire __A17_2__CCH10;
    wire __A17_2__RCH10_n;
    wire __A17_2__WCH10_n;
    wire __A17_NET_176;
    wire __A17_NET_176_U17019_10;
    wire __A17_NET_176_U17019_8;
    wire __A17_NET_177;
    wire __A17_NET_178;
    wire __A17_NET_179;
    wire __A17_NET_180;
    wire __A17_NET_181;
    wire __A17_NET_182;
    wire __A17_NET_183;
    wire __A17_NET_183_U17019_12;
    wire __A17_NET_183_U17027_2;
    wire __A17_NET_184;
    wire __A17_NET_185;
    wire __A17_NET_186;
    wire __A17_NET_187;
    wire __A17_NET_188;
    wire __A17_NET_189;
    wire __A17_NET_190;
    wire __A17_NET_191;
    wire __A17_NET_192;
    wire __A17_NET_193;
    wire __A17_NET_194;
    wire __A17_NET_195;
    wire __A17_NET_196;
    wire __A17_NET_197;
    wire __A17_NET_198;
    wire __A17_NET_199;
    wire __A17_NET_200;
    wire __A17_NET_201;
    wire __A17_NET_202;
    wire __A17_NET_203;
    wire __A17_NET_204;
    wire __A17_NET_205;
    wire __A17_NET_206;
    wire __A17_NET_207;
    wire __A17_NET_208;
    wire __A17_NET_209;
    wire __A17_NET_210;
    wire __A17_NET_211;
    wire __A17_NET_212;
    wire __A17_NET_213;
    wire __A17_NET_214;
    wire __A17_NET_215;
    wire __A17_NET_216;
    wire __A17_NET_217;
    wire __A17_NET_218;
    wire __A17_NET_219;
    wire __A17_NET_220;
    wire __A17_NET_220_U17027_4;
    wire __A17_NET_220_U17027_6;
    wire __A17_NET_220_U17027_8;
    wire __A17_NET_221;
    wire __A17_NET_222;
    wire __A17_NET_225;
    wire __A17_NET_226;
    wire __A17_NET_227;
    wire __A17_NET_228;
    wire __A17_NET_229;
    wire __A17_NET_230;
    wire __A17_NET_231;
    wire __A17_NET_232;
    wire __A17_NET_233;
    wire __A17_NET_234;
    wire __A17_NET_235;
    wire __A17_NET_236;
    wire __A17_NET_237;
    wire __A17_NET_238;
    wire __A17_NET_239;
    wire __A17_NET_240;
    wire __A17_NET_241;
    wire __A17_NET_242;
    wire __A17_NET_243;
    wire __A17_NET_244;
    wire __A17_NET_245;
    wire __A17_NET_246;
    wire __A17_NET_247;
    wire __A17_NET_248;
    wire __A17_NET_249;
    wire __A17_NET_250;
    wire __A17_NET_251;
    wire __A17_NET_252;
    wire __A17_NET_253;
    wire __A17_NET_254;
    wire __A17_NET_255;
    wire __A17_NET_256;
    wire __A17_NET_257;
    wire __A17_NET_258;
    wire __A17_NET_259;
    wire __A17_NET_260;
    wire __A17_NET_261;
    wire __A17_NET_262;
    wire __A17_NET_263;
    wire __A17_NET_264;
    wire __A17_NET_265;
    wire __A17_NET_266;
    wire __A17_NET_267;
    wire __A17_NET_269;
    wire __A17_NET_270;
    wire __A17_NET_271;
    wire __A17_NET_272;
    wire __A17_NET_273;
    wire __A17_NET_274;
    wire __A17_NET_275;
    wire __A17_NET_276;
    wire __A17_NET_277;
    wire __A17_NET_278;
    wire __A17_NET_279;
    wire __A17_NET_280;
    wire __A17_NET_281;
    wire __A17_NET_282;
    wire __A17_NET_283;
    wire __A17_NET_284;
    wire __A17_NET_285;
    wire __A17_NET_286;
    wire __A17_NET_287;
    wire __A17_NET_288;
    wire __A17_NET_289;
    wire __A17_NET_290;
    wire __A17_NET_291;
    wire __A17_NET_292;
    wire __A17_NET_293;
    wire __A17_NET_294;
    wire __A17_NET_295;
    wire __A17_NET_296;
    wire __A17_NET_297;
    wire __A17_NET_298;
    wire __A17_NET_299;
    wire __A17_NET_300;
    wire __A17_NET_301;
    wire __A17_NET_302;
    wire __A17_NET_303;
    wire __A17_NET_304;
    wire __A17_NET_305;
    wire __A17_NET_306;
    wire __A17_NET_307;
    wire __A17_NET_308;
    wire __A17_NET_309;
    wire __A17_NET_310;
    wire __A17_NET_311;
    wire __A17_NET_312;
    wire __A17_NET_313;
    wire __A17_NET_314;
    wire __A17_NET_315;
    wire __A17_NET_316;
    wire __A17_NET_318;
    wire __A17_NET_319;
    wire __A17_NET_320;
    wire __A17_NET_321;
    wire __A17_NET_322;
    wire __A17_NET_323;
    wire __A17_NET_324;
    wire __A17_NET_325;
    wire __A17_NET_326;
    wire __A17_NET_327;
    wire __A17_NET_328;
    wire __A17_NET_329;
    wire __A17_NET_330;
    wire __A17_NET_331;
    wire __A17_NET_332;
    wire __A17_NET_333;
    wire __A17_NET_334;
    wire __A17_NET_335;
    wire __A17_NET_336;
    wire __A17_NET_337;
    wire __A17_NET_338;
    wire __A17_NET_339;
    wire __A17_NET_340;
    wire __A17_NET_341;
    wire __A17_NET_342;
    wire __A17_NET_343;
    wire __A17_NET_344;
    wire __A17_NET_346;
    wire __A17_NET_347;
    wire __A17_NET_348;
    wire __A17_NET_349;
    wire __A17_NET_350;
    wire __A17_NET_351;
    wire __A17_NET_352;
    wire __A17_NET_354;
    wire __A17_NET_355;
    wire __A17_NET_356;
    wire __A18_1__F08B_n;
    wire __A18_1__F09A_n;
    wire __A18_1__F09D;
    wire __A18_1__F17A_n;
    wire __A18_1__F17B_n;
    wire __A18_1__RCH15_n;
    wire __A18_1__RCH16_n;
    wire __A18_1__STNDBY;
    wire __A18_2__ACTV_n;
    wire __A18_2__ADVCNT;
    wire __A18_2__CNTOF9;
    wire __A18_2__CNTOF9_U18007_10;
    wire __A18_2__CNTOF9_U18007_12;
    wire __A18_2__F10AS0;
    wire __A18_2__HERB;
    wire __A18_2__LRRANG;
    wire __A18_2__LRSYNC;
    wire __A18_2__LRXVEL;
    wire __A18_2__LRYVEL;
    wire __A18_2__LRZVEL;
    wire __A18_2__RRRANG;
    wire __A18_2__RRRARA;
    wire __A18_2__RRSYNC;
    wire __A18_NET_100;
    wire __A18_NET_101;
    wire __A18_NET_102;
    wire __A18_NET_103;
    wire __A18_NET_104;
    wire __A18_NET_105;
    wire __A18_NET_106;
    wire __A18_NET_107;
    wire __A18_NET_108;
    wire __A18_NET_109;
    wire __A18_NET_110;
    wire __A18_NET_111;
    wire __A18_NET_112;
    wire __A18_NET_113;
    wire __A18_NET_114;
    wire __A18_NET_116;
    wire __A18_NET_116_U18007_2;
    wire __A18_NET_116_U18007_4;
    wire __A18_NET_117;
    wire __A18_NET_118;
    wire __A18_NET_119;
    wire __A18_NET_120;
    wire __A18_NET_121;
    wire __A18_NET_122;
    wire __A18_NET_123;
    wire __A18_NET_124;
    wire __A18_NET_125;
    wire __A18_NET_126;
    wire __A18_NET_127;
    wire __A18_NET_128;
    wire __A18_NET_129;
    wire __A18_NET_130;
    wire __A18_NET_131;
    wire __A18_NET_132;
    wire __A18_NET_133;
    wire __A18_NET_134;
    wire __A18_NET_135;
    wire __A18_NET_136;
    wire __A18_NET_137;
    wire __A18_NET_138;
    wire __A18_NET_139;
    wire __A18_NET_140;
    wire __A18_NET_141;
    wire __A18_NET_142;
    wire __A18_NET_143;
    wire __A18_NET_144;
    wire __A18_NET_145;
    wire __A18_NET_146;
    wire __A18_NET_147;
    wire __A18_NET_149;
    wire __A18_NET_150;
    wire __A18_NET_151;
    wire __A18_NET_155;
    wire __A18_NET_156;
    wire __A18_NET_157;
    wire __A18_NET_158;
    wire __A18_NET_159;
    wire __A18_NET_160;
    wire __A18_NET_161;
    wire __A18_NET_162;
    wire __A18_NET_163;
    wire __A18_NET_164;
    wire __A18_NET_165;
    wire __A18_NET_166;
    wire __A18_NET_167;
    wire __A18_NET_168;
    wire __A18_NET_169;
    wire __A18_NET_170;
    wire __A18_NET_171;
    wire __A18_NET_172;
    wire __A18_NET_173;
    wire __A18_NET_174;
    wire __A18_NET_178;
    wire __A18_NET_179;
    wire __A18_NET_180;
    wire __A18_NET_181;
    wire __A18_NET_182;
    wire __A18_NET_184;
    wire __A18_NET_187;
    wire __A18_NET_188;
    wire __A18_NET_189;
    wire __A18_NET_192;
    wire __A18_NET_193;
    wire __A18_NET_194;
    wire __A18_NET_195;
    wire __A18_NET_196;
    wire __A18_NET_197;
    wire __A18_NET_198;
    wire __A18_NET_199;
    wire __A18_NET_200;
    wire __A18_NET_201;
    wire __A18_NET_202;
    wire __A18_NET_203;
    wire __A18_NET_204;
    wire __A18_NET_205;
    wire __A18_NET_206;
    wire __A18_NET_207;
    wire __A18_NET_208;
    wire __A18_NET_209;
    wire __A18_NET_210;
    wire __A18_NET_211;
    wire __A18_NET_212;
    wire __A18_NET_213;
    wire __A18_NET_214;
    wire __A18_NET_216;
    wire __A18_NET_217;
    wire __A18_NET_218;
    wire __A18_NET_219;
    wire __A18_NET_220;
    wire __A18_NET_221;
    wire __A18_NET_222;
    wire __A18_NET_223;
    wire __A18_NET_224;
    wire __A18_NET_225;
    wire __A18_NET_226;
    wire __A18_NET_227;
    wire __A18_NET_228;
    wire __A18_NET_229;
    wire __A18_NET_230;
    wire __A18_NET_231;
    wire __A18_NET_232;
    wire __A18_NET_233;
    wire __A18_NET_234;
    wire __A18_NET_235;
    wire __A18_NET_238;
    wire __A18_NET_241;
    wire __A18_NET_242;
    wire __A18_NET_247;
    wire __A18_NET_248;
    wire __A18_NET_249;
    wire __A18_NET_250;
    wire __A18_NET_251;
    wire __A18_NET_253;
    wire __A18_NET_254;
    wire __A18_NET_256;
    wire __A18_NET_257;
    wire __A18_NET_258;
    wire __A18_NET_259;
    wire __A18_NET_260;
    wire __A18_NET_261;
    wire __A18_NET_262;
    wire __A18_NET_263;
    wire __A18_NET_264;
    wire __A18_NET_265;
    wire __A18_NET_266;
    wire __A18_NET_267;
    wire __A18_NET_268;
    wire __A18_NET_269;
    wire __A18_NET_270;
    wire __A18_NET_272;
    wire __A18_NET_273;
    wire __A18_NET_274;
    wire __A18_NET_275;
    wire __A18_NET_276;
    wire __A18_NET_93;
    wire __A18_NET_94;
    wire __A18_NET_95;
    wire __A18_NET_96;
    wire __A18_NET_97;
    wire __A18_NET_98;
    wire __A18_NET_99;
    wire __A18_NET_99_U18007_6;
    wire __A18_NET_99_U18007_8;
    wire __A19_1__ALRT0;
    wire __A19_1__ALRT1;
    wire __A19_1__ALT0;
    wire __A19_1__ALT1;
    wire __A19_1__ALTSNC;
    wire __A19_1__BLKUPL;
    wire __A19_1__C45R_n;
    wire __A19_1__EMSm;
    wire __A19_1__EMSp;
    wire __A19_1__F5ASB0;
    wire __A19_1__F5BSB2;
    wire __A19_1__OTLNK0;
    wire __A19_1__OTLNK1;
    wire __A19_1__SH3MS_n;
    wire __A19_1__THRSTm;
    wire __A19_1__THRSTp;
    wire __A19_1__UPL0_n;
    wire __A19_1__UPL1_n;
    wire __A19_1__XLNK0_n;
    wire __A19_1__XLNK1_n;
    wire __A19_2__CNTRSB_n;
    wire __A19_2__F06B_n;
    wire __A19_2__F07C_n;
    wire __A19_2__F07D_n;
    wire __A19_2__F10B_n;
    wire __A19_2__F7CSB1_n;
    wire __A19_2__FF1109_n;
    wire __A19_2__FF1110_n;
    wire __A19_2__FF1111_n;
    wire __A19_2__FF1112_n;
    wire __A19_2__GYENAB;
    wire __A19_2__GYRRST;
    wire __A19_2__GYRSET;
    wire __A19_2__GYXM;
    wire __A19_2__GYXP;
    wire __A19_2__GYYM;
    wire __A19_2__GYYP;
    wire __A19_2__GYZM;
    wire __A19_2__GYZP;
    wire __A19_2__O44;
    wire __A19_2__OT1110;
    wire __A19_2__OT1111;
    wire __A19_2__OT1112;
    wire __A19_2__RHCGO;
    wire __A19_NET_159;
    wire __A19_NET_161;
    wire __A19_NET_162;
    wire __A19_NET_163;
    wire __A19_NET_164;
    wire __A19_NET_165;
    wire __A19_NET_166;
    wire __A19_NET_167;
    wire __A19_NET_168;
    wire __A19_NET_169;
    wire __A19_NET_170;
    wire __A19_NET_171;
    wire __A19_NET_172;
    wire __A19_NET_173;
    wire __A19_NET_176;
    wire __A19_NET_177;
    wire __A19_NET_178;
    wire __A19_NET_179;
    wire __A19_NET_180;
    wire __A19_NET_181;
    wire __A19_NET_182;
    wire __A19_NET_184;
    wire __A19_NET_185;
    wire __A19_NET_186;
    wire __A19_NET_187;
    wire __A19_NET_188;
    wire __A19_NET_189;
    wire __A19_NET_190;
    wire __A19_NET_192;
    wire __A19_NET_193;
    wire __A19_NET_194;
    wire __A19_NET_195;
    wire __A19_NET_196;
    wire __A19_NET_197;
    wire __A19_NET_198;
    wire __A19_NET_199;
    wire __A19_NET_200;
    wire __A19_NET_201;
    wire __A19_NET_202;
    wire __A19_NET_203;
    wire __A19_NET_204;
    wire __A19_NET_205;
    wire __A19_NET_206;
    wire __A19_NET_207;
    wire __A19_NET_208;
    wire __A19_NET_209;
    wire __A19_NET_210;
    wire __A19_NET_211;
    wire __A19_NET_212;
    wire __A19_NET_213;
    wire __A19_NET_214;
    wire __A19_NET_215;
    wire __A19_NET_216;
    wire __A19_NET_217;
    wire __A19_NET_218;
    wire __A19_NET_219;
    wire __A19_NET_220;
    wire __A19_NET_221;
    wire __A19_NET_222;
    wire __A19_NET_223;
    wire __A19_NET_224;
    wire __A19_NET_225;
    wire __A19_NET_226;
    wire __A19_NET_227;
    wire __A19_NET_228;
    wire __A19_NET_229;
    wire __A19_NET_230;
    wire __A19_NET_231;
    wire __A19_NET_232;
    wire __A19_NET_234;
    wire __A19_NET_235;
    wire __A19_NET_236;
    wire __A19_NET_238;
    wire __A19_NET_241;
    wire __A19_NET_242;
    wire __A19_NET_243;
    wire __A19_NET_244;
    wire __A19_NET_245;
    wire __A19_NET_246;
    wire __A19_NET_247;
    wire __A19_NET_248;
    wire __A19_NET_249;
    wire __A19_NET_250;
    wire __A19_NET_251;
    wire __A19_NET_252;
    wire __A19_NET_253;
    wire __A19_NET_254;
    wire __A19_NET_255;
    wire __A19_NET_256;
    wire __A19_NET_257;
    wire __A19_NET_258;
    wire __A19_NET_259;
    wire __A19_NET_260;
    wire __A19_NET_261;
    wire __A19_NET_262;
    wire __A19_NET_263;
    wire __A19_NET_264;
    wire __A19_NET_265;
    wire __A19_NET_266;
    wire __A19_NET_267;
    wire __A19_NET_268;
    wire __A19_NET_269;
    wire __A19_NET_270;
    wire __A19_NET_271;
    wire __A19_NET_272;
    wire __A19_NET_273;
    wire __A19_NET_274;
    wire __A19_NET_275;
    wire __A19_NET_276;
    wire __A19_NET_277;
    wire __A19_NET_278;
    wire __A19_NET_279;
    wire __A19_NET_280;
    wire __A19_NET_281;
    wire __A19_NET_282;
    wire __A19_NET_283;
    wire __A19_NET_284;
    wire __A19_NET_285;
    wire __A19_NET_286;
    wire __A19_NET_287;
    wire __A19_NET_289;
    wire __A19_NET_290;
    wire __A19_NET_291;
    wire __A19_NET_292;
    wire __A19_NET_293;
    wire __A19_NET_299;
    wire __A19_NET_300;
    wire __A19_NET_301;
    wire __A19_NET_302;
    wire __A19_NET_303;
    wire __A19_NET_304;
    wire __A19_NET_305;
    wire __A19_NET_306;
    wire __A19_NET_307;
    wire __A19_NET_308;
    wire __A19_NET_309;
    wire __A19_NET_310;
    wire __A19_NET_311;
    wire __A19_NET_312;
    wire __A19_NET_314;
    wire __A19_NET_315;
    wire __A19_NET_316;
    wire __A19_NET_317;
    wire __A19_NET_318;
    wire __A19_NET_319;
    wire __A19_NET_320;
    wire __A19_NET_321;
    wire __A19_NET_322;
    wire __A19_NET_323;
    wire __A19_NET_325;
    wire __A19_NET_326;
    wire __A19_NET_328;
    wire __A19_NET_329;
    wire __A19_NET_330;
    wire __A20_1__C10R;
    wire __A20_1__C1R;
    wire __A20_1__C2R;
    wire __A20_1__C3R;
    wire __A20_1__C4R;
    wire __A20_1__C5R;
    wire __A20_1__C6R;
    wire __A20_1__C7R;
    wire __A20_1__C8R;
    wire __A20_1__C9R;
    wire __A20_2__C10R;
    wire __A20_2__C1R;
    wire __A20_2__C2R;
    wire __A20_2__C3R;
    wire __A20_2__C4R;
    wire __A20_2__C5R;
    wire __A20_2__C6R;
    wire __A20_2__C7R;
    wire __A20_2__C8R;
    wire __A20_2__C9R;
    wire __A20_NET_100;
    wire __A20_NET_101;
    wire __A20_NET_102;
    wire __A20_NET_103;
    wire __A20_NET_104;
    wire __A20_NET_105;
    wire __A20_NET_107;
    wire __A20_NET_108;
    wire __A20_NET_109;
    wire __A20_NET_110;
    wire __A20_NET_111;
    wire __A20_NET_112;
    wire __A20_NET_113;
    wire __A20_NET_115;
    wire __A20_NET_120;
    wire __A20_NET_121;
    wire __A20_NET_122;
    wire __A20_NET_123;
    wire __A20_NET_124;
    wire __A20_NET_125;
    wire __A20_NET_127;
    wire __A20_NET_128;
    wire __A20_NET_129;
    wire __A20_NET_130;
    wire __A20_NET_131;
    wire __A20_NET_132;
    wire __A20_NET_134;
    wire __A20_NET_135;
    wire __A20_NET_136;
    wire __A20_NET_137;
    wire __A20_NET_138;
    wire __A20_NET_139;
    wire __A20_NET_140;
    wire __A20_NET_142;
    wire __A20_NET_143;
    wire __A20_NET_144;
    wire __A20_NET_145;
    wire __A20_NET_146;
    wire __A20_NET_147;
    wire __A20_NET_148;
    wire __A20_NET_150;
    wire __A20_NET_151;
    wire __A20_NET_152;
    wire __A20_NET_153;
    wire __A20_NET_155;
    wire __A20_NET_156;
    wire __A20_NET_157;
    wire __A20_NET_158;
    wire __A20_NET_160;
    wire __A20_NET_161;
    wire __A20_NET_165;
    wire __A20_NET_166;
    wire __A20_NET_167;
    wire __A20_NET_168;
    wire __A20_NET_170;
    wire __A20_NET_171;
    wire __A20_NET_172;
    wire __A20_NET_173;
    wire __A20_NET_175;
    wire __A20_NET_176;
    wire __A20_NET_177;
    wire __A20_NET_178;
    wire __A20_NET_179;
    wire __A20_NET_180;
    wire __A20_NET_181;
    wire __A20_NET_182;
    wire __A20_NET_184;
    wire __A20_NET_185;
    wire __A20_NET_186;
    wire __A20_NET_187;
    wire __A20_NET_188;
    wire __A20_NET_189;
    wire __A20_NET_190;
    wire __A20_NET_191;
    wire __A20_NET_192;
    wire __A20_NET_194;
    wire __A20_NET_195;
    wire __A20_NET_196;
    wire __A20_NET_197;
    wire __A20_NET_198;
    wire __A20_NET_199;
    wire __A20_NET_200;
    wire __A20_NET_201;
    wire __A20_NET_203;
    wire __A20_NET_208;
    wire __A20_NET_209;
    wire __A20_NET_210;
    wire __A20_NET_211;
    wire __A20_NET_212;
    wire __A20_NET_213;
    wire __A20_NET_215;
    wire __A20_NET_216;
    wire __A20_NET_217;
    wire __A20_NET_218;
    wire __A20_NET_219;
    wire __A20_NET_220;
    wire __A20_NET_222;
    wire __A20_NET_223;
    wire __A20_NET_224;
    wire __A20_NET_225;
    wire __A20_NET_226;
    wire __A20_NET_227;
    wire __A20_NET_228;
    wire __A20_NET_230;
    wire __A20_NET_231;
    wire __A20_NET_232;
    wire __A20_NET_233;
    wire __A20_NET_234;
    wire __A20_NET_235;
    wire __A20_NET_236;
    wire __A20_NET_237;
    wire __A20_NET_239;
    wire __A20_NET_240;
    wire __A20_NET_241;
    wire __A20_NET_243;
    wire __A20_NET_244;
    wire __A20_NET_245;
    wire __A20_NET_246;
    wire __A20_NET_247;
    wire __A20_NET_250;
    wire __A20_NET_251;
    wire __A20_NET_254;
    wire __A20_NET_255;
    wire __A20_NET_256;
    wire __A20_NET_258;
    wire __A20_NET_259;
    wire __A20_NET_260;
    wire __A20_NET_261;
    wire __A20_NET_263;
    wire __A20_NET_264;
    wire __A20_NET_265;
    wire __A20_NET_90;
    wire __A20_NET_91;
    wire __A20_NET_92;
    wire __A20_NET_93;
    wire __A20_NET_94;
    wire __A20_NET_96;
    wire __A20_NET_97;
    wire __A20_NET_98;
    wire __A20_NET_99;
    wire __A21_1__30SUM;
    wire __A21_1__32004K;
    wire __A21_1__32004K_U21010_2;
    wire __A21_1__32004K_U21010_4;
    wire __A21_1__50SUM;
    wire __A21_1__C42A;
    wire __A21_1__C42M;
    wire __A21_1__C42P;
    wire __A21_1__C43A;
    wire __A21_1__C43M;
    wire __A21_1__C43P;
    wire __A21_1__C44A;
    wire __A21_1__C44M;
    wire __A21_1__C44P;
    wire __A21_1__C45A;
    wire __A21_1__C45M;
    wire __A21_1__C45P;
    wire __A21_1__C46A;
    wire __A21_1__C46M;
    wire __A21_1__C46P;
    wire __A21_1__C47A;
    wire __A21_1__C56A;
    wire __A21_1__C57A;
    wire __A21_1__C60A;
    wire __A21_1__DINCNC_n;
    wire __A21_1__MCDU_n;
    wire __A21_1__MINC_n;
    wire __A21_1__PCDU_n;
    wire __A21_1__PINC_n;
    wire __A21_1__RSCT_n;
    wire __A21_1__SHANC;
    wire __A21_1__SHINC;
    wire __A21_3__C42R;
    wire __A21_3__C43R;
    wire __A21_3__C44R;
    wire __A21_3__C46R;
    wire __A21_3__C47R;
    wire __A21_3__C56R;
    wire __A21_3__C57R;
    wire __A21_3__C60R;
    wire __A21_3__CG15;
    wire __A21_3__CG16;
    wire __A21_NET_133;
    wire __A21_NET_134;
    wire __A21_NET_136;
    wire __A21_NET_140;
    wire __A21_NET_141;
    wire __A21_NET_141_U21023_2;
    wire __A21_NET_141_U21023_4;
    wire __A21_NET_141_U21023_6;
    wire __A21_NET_142;
    wire __A21_NET_143;
    wire __A21_NET_144;
    wire __A21_NET_145;
    wire __A21_NET_145_U21023_10;
    wire __A21_NET_145_U21023_8;
    wire __A21_NET_146;
    wire __A21_NET_146_U21010_10;
    wire __A21_NET_146_U21010_12;
    wire __A21_NET_147;
    wire __A21_NET_147_U21006_10;
    wire __A21_NET_147_U21006_12;
    wire __A21_NET_147_U21006_6;
    wire __A21_NET_147_U21006_8;
    wire __A21_NET_148;
    wire __A21_NET_149;
    wire __A21_NET_151;
    wire __A21_NET_152;
    wire __A21_NET_152_U21002_2;
    wire __A21_NET_152_U21002_4;
    wire __A21_NET_152_U21002_6;
    wire __A21_NET_152_U21002_8;
    wire __A21_NET_153;
    wire __A21_NET_153_U21002_10;
    wire __A21_NET_153_U21002_12;
    wire __A21_NET_153_U21006_2;
    wire __A21_NET_153_U21006_4;
    wire __A21_NET_154;
    wire __A21_NET_156;
    wire __A21_NET_157;
    wire __A21_NET_159;
    wire __A21_NET_159_U21023_12;
    wire __A21_NET_159_U21027_2;
    wire __A21_NET_160;
    wire __A21_NET_161;
    wire __A21_NET_162;
    wire __A21_NET_162_U21027_4;
    wire __A21_NET_162_U21027_6;
    wire __A21_NET_163;
    wire __A21_NET_164;
    wire __A21_NET_165;
    wire __A21_NET_166;
    wire __A21_NET_168;
    wire __A21_NET_172;
    wire __A21_NET_173;
    wire __A21_NET_173_U21010_6;
    wire __A21_NET_173_U21010_8;
    wire __A21_NET_174;
    wire __A21_NET_178;
    wire __A21_NET_179;
    wire __A21_NET_184;
    wire __A21_NET_185;
    wire __A21_NET_187;
    wire __A21_NET_187_U21014_2;
    wire __A21_NET_187_U21014_4;
    wire __A21_NET_187_U21014_6;
    wire __A21_NET_188;
    wire __A21_NET_193;
    wire __A21_NET_194;
    wire __A21_NET_199;
    wire __A21_NET_200;
    wire __A21_NET_203;
    wire __A21_NET_204;
    wire __A21_NET_205;
    wire __A21_NET_212;
    wire __A21_NET_215;
    wire __A21_NET_216;
    wire __A21_NET_219;
    wire __A21_NET_224;
    wire __A21_NET_225;
    wire __A21_NET_226;
    wire __A21_NET_227;
    wire __A21_NET_228;
    wire __A21_NET_229;
    wire __A21_NET_229_U21014_10;
    wire __A21_NET_229_U21014_12;
    wire __A21_NET_229_U21014_8;
    wire __A21_NET_232;
    wire __A21_NET_233;
    wire __A21_NET_234;
    wire __A21_NET_235;
    wire __A21_NET_236;
    wire __A21_NET_237;
    wire __A21_NET_238;
    wire __A21_NET_239;
    wire __A21_NET_240;
    wire __A21_NET_241;
    wire __A21_NET_242;
    wire __A21_NET_243;
    wire __A21_NET_244;
    wire __A21_NET_245;
    wire __A21_NET_246;
    wire __A21_NET_247;
    wire __A21_NET_248;
    wire __A21_NET_249;
    wire __A21_NET_250;
    wire __A21_NET_251;
    wire __A21_NET_252;
    wire __A21_NET_253;
    wire __A21_NET_254;
    wire __A21_NET_255;
    wire __A21_NET_256;
    wire __A21_NET_257;
    wire __A21_NET_258;
    wire __A21_NET_259;
    wire __A21_NET_260;
    wire __A21_NET_261;
    wire __A21_NET_262;
    wire __A21_NET_263;
    wire __A21_NET_264;
    wire __A21_NET_265;
    wire __A21_NET_266;
    wire __A21_NET_267;
    wire __A21_NET_268;
    wire __A21_NET_269;
    wire __A21_NET_271;
    wire __A21_NET_272;
    wire __A21_NET_273;
    wire __A21_NET_274;
    wire __A21_NET_275;
    wire __A21_NET_276;
    wire __A21_NET_277;
    wire __A21_NET_278;
    wire __A21_NET_279;
    wire __A21_NET_280;
    wire __A21_NET_281;
    wire __A21_NET_282;
    wire __A21_NET_283;
    wire __A21_NET_284;
    wire __A21_NET_285;
    wire __A21_NET_286;
    wire __A21_NET_287;
    wire __A21_NET_288;
    wire __A21_NET_289;
    wire __A21_NET_290;
    wire __A21_NET_292;
    wire __A21_NET_300;
    wire __A21_NET_301;
    wire __A21_NET_302;
    wire __A21_NET_304;
    wire __A21_NET_305;
    wire __A21_NET_306;
    wire __A21_NET_307;
    wire __A21_NET_308;
    wire __A21_NET_71;
    wire __A22_1__16CNT;
    wire __A22_1__1CNT;
    wire __A22_1__32CNT;
    wire __A22_1__ADVCTR;
    wire __A22_1__BSYNC_n;
    wire __A22_1__DATA_n;
    wire __A22_1__DATA_n_U22028_10;
    wire __A22_1__DATA_n_U22028_12;
    wire __A22_1__DATA_n_U22028_2;
    wire __A22_1__DATA_n_U22028_4;
    wire __A22_1__DATA_n_U22028_6;
    wire __A22_1__DATA_n_U22028_8;
    wire __A22_1__DATA_n_U22057_2;
    wire __A22_1__DATA_n_U22057_4;
    wire __A22_1__DATA_n_U22057_6;
    wire __A22_1__DKCTR1;
    wire __A22_1__DKCTR1_n;
    wire __A22_1__DKCTR2;
    wire __A22_1__DKCTR2_n;
    wire __A22_1__DKCTR3;
    wire __A22_1__DKCTR3_n;
    wire __A22_1__DKCTR4;
    wire __A22_1__DKCTR4_n;
    wire __A22_1__DKCTR5;
    wire __A22_1__DKCTR5_n;
    wire __A22_1__DKDATB;
    wire __A22_1__DKDAT_n;
    wire __A22_1__DLKCLR;
    wire __A22_1__DLKRPT;
    wire __A22_1__END;
    wire __A22_1__HIGH0_n;
    wire __A22_1__HIGH1_n;
    wire __A22_1__HIGH2_n;
    wire __A22_1__HIGH3_n;
    wire __A22_1__LOW0_n;
    wire __A22_1__LOW1_n;
    wire __A22_1__LOW2_n;
    wire __A22_1__LOW3_n;
    wire __A22_1__LOW4_n;
    wire __A22_1__LOW5_n;
    wire __A22_1__LOW6_n;
    wire __A22_1__LOW7_n;
    wire __A22_1__ORDRBT;
    wire __A22_1__RDOUT_n;
    wire __A22_1__WDORDR;
    wire __A22_1__WRD1B1;
    wire __A22_1__WRD1BP;
    wire __A22_1__WRD2B2;
    wire __A22_1__WRD2B3;
    wire __A22_NET_100;
    wire __A22_NET_102;
    wire __A22_NET_103;
    wire __A22_NET_104;
    wire __A22_NET_105;
    wire __A22_NET_107;
    wire __A22_NET_108;
    wire __A22_NET_109;
    wire __A22_NET_111;
    wire __A22_NET_112;
    wire __A22_NET_116;
    wire __A22_NET_117;
    wire __A22_NET_118;
    wire __A22_NET_119;
    wire __A22_NET_120;
    wire __A22_NET_121;
    wire __A22_NET_122;
    wire __A22_NET_123;
    wire __A22_NET_124;
    wire __A22_NET_125;
    wire __A22_NET_127;
    wire __A22_NET_128;
    wire __A22_NET_129;
    wire __A22_NET_130;
    wire __A22_NET_131;
    wire __A22_NET_132;
    wire __A22_NET_133;
    wire __A22_NET_135;
    wire __A22_NET_136;
    wire __A22_NET_137;
    wire __A22_NET_138;
    wire __A22_NET_139;
    wire __A22_NET_140;
    wire __A22_NET_141;
    wire __A22_NET_142;
    wire __A22_NET_143;
    wire __A22_NET_144;
    wire __A22_NET_145;
    wire __A22_NET_146;
    wire __A22_NET_147;
    wire __A22_NET_148;
    wire __A22_NET_149;
    wire __A22_NET_150;
    wire __A22_NET_151;
    wire __A22_NET_152;
    wire __A22_NET_153;
    wire __A22_NET_154;
    wire __A22_NET_155;
    wire __A22_NET_156;
    wire __A22_NET_157;
    wire __A22_NET_158;
    wire __A22_NET_159;
    wire __A22_NET_160;
    wire __A22_NET_161;
    wire __A22_NET_162;
    wire __A22_NET_163;
    wire __A22_NET_164;
    wire __A22_NET_167;
    wire __A22_NET_168;
    wire __A22_NET_169;
    wire __A22_NET_170;
    wire __A22_NET_171;
    wire __A22_NET_172;
    wire __A22_NET_173;
    wire __A22_NET_174;
    wire __A22_NET_175;
    wire __A22_NET_176;
    wire __A22_NET_177;
    wire __A22_NET_180;
    wire __A22_NET_181;
    wire __A22_NET_182;
    wire __A22_NET_183;
    wire __A22_NET_184;
    wire __A22_NET_185;
    wire __A22_NET_186;
    wire __A22_NET_187;
    wire __A22_NET_188;
    wire __A22_NET_189;
    wire __A22_NET_190;
    wire __A22_NET_191;
    wire __A22_NET_192;
    wire __A22_NET_193;
    wire __A22_NET_194;
    wire __A22_NET_195;
    wire __A22_NET_196;
    wire __A22_NET_197;
    wire __A22_NET_198;
    wire __A22_NET_199;
    wire __A22_NET_200;
    wire __A22_NET_201;
    wire __A22_NET_202;
    wire __A22_NET_203;
    wire __A22_NET_204;
    wire __A22_NET_205;
    wire __A22_NET_206;
    wire __A22_NET_207;
    wire __A22_NET_208;
    wire __A22_NET_209;
    wire __A22_NET_210;
    wire __A22_NET_211;
    wire __A22_NET_213;
    wire __A22_NET_214;
    wire __A22_NET_215;
    wire __A22_NET_217;
    wire __A22_NET_218;
    wire __A22_NET_219;
    wire __A22_NET_220;
    wire __A22_NET_221;
    wire __A22_NET_222;
    wire __A22_NET_223;
    wire __A22_NET_224;
    wire __A22_NET_225;
    wire __A22_NET_226;
    wire __A22_NET_227;
    wire __A22_NET_228;
    wire __A22_NET_229;
    wire __A22_NET_230;
    wire __A22_NET_231;
    wire __A22_NET_232;
    wire __A22_NET_233;
    wire __A22_NET_234;
    wire __A22_NET_235;
    wire __A22_NET_236;
    wire __A22_NET_237;
    wire __A22_NET_238;
    wire __A22_NET_239;
    wire __A22_NET_240;
    wire __A22_NET_241;
    wire __A22_NET_242;
    wire __A22_NET_243;
    wire __A22_NET_244;
    wire __A22_NET_245;
    wire __A22_NET_246;
    wire __A22_NET_247;
    wire __A22_NET_248;
    wire __A22_NET_251;
    wire __A22_NET_252;
    wire __A22_NET_253;
    wire __A22_NET_254;
    wire __A22_NET_255;
    wire __A22_NET_256;
    wire __A22_NET_257;
    wire __A22_NET_258;
    wire __A22_NET_259;
    wire __A22_NET_261;
    wire __A22_NET_262;
    wire __A22_NET_263;
    wire __A22_NET_265;
    wire __A22_NET_266;
    wire __A22_NET_267;
    wire __A22_NET_268;
    wire __A22_NET_269;
    wire __A22_NET_270;
    wire __A22_NET_271;
    wire __A22_NET_272;
    wire __A22_NET_273;
    wire __A22_NET_274;
    wire __A22_NET_275;
    wire __A22_NET_276;
    wire __A22_NET_279;
    wire __A22_NET_280;
    wire __A22_NET_281;
    wire __A22_NET_282;
    wire __A22_NET_283;
    wire __A22_NET_284;
    wire __A22_NET_285;
    wire __A22_NET_286;
    wire __A22_NET_287;
    wire __A22_NET_58;
    wire __A22_NET_60;
    wire __A22_NET_61;
    wire __A22_NET_64;
    wire __A22_NET_66;
    wire __A22_NET_67;
    wire __A22_NET_68;
    wire __A22_NET_69;
    wire __A22_NET_71;
    wire __A22_NET_74;
    wire __A22_NET_75;
    wire __A22_NET_78;
    wire __A22_NET_79;
    wire __A22_NET_80;
    wire __A22_NET_81;
    wire __A22_NET_82;
    wire __A22_NET_83;
    wire __A22_NET_84;
    wire __A22_NET_85;
    wire __A22_NET_86;
    wire __A22_NET_87;
    wire __A22_NET_88;
    wire __A22_NET_89;
    wire __A22_NET_90;
    wire __A22_NET_91;
    wire __A22_NET_92;
    wire __A22_NET_95;
    wire __A22_NET_96;
    wire __A23_1__BOTHX;
    wire __A23_1__BOTHY;
    wire __A23_1__BOTHZ;
    wire __A23_1__F18AX;
    wire __A23_1__F18A_n;
    wire __A23_1__F18B_n;
    wire __A23_1__MISSX;
    wire __A23_1__MISSY;
    wire __A23_1__MISSZ;
    wire __A23_1__NOXM;
    wire __A23_1__NOXP;
    wire __A23_1__NOYM;
    wire __A23_1__NOYP;
    wire __A23_1__NOZM;
    wire __A23_1__NOZP;
    wire __A23_1__P04A;
    wire __A23_1__PIPAXm_n;
    wire __A23_1__PIPAXp_n;
    wire __A23_1__PIPAYm_n;
    wire __A23_1__PIPAYp_n;
    wire __A23_1__PIPAZm_n;
    wire __A23_1__PIPAZp_n;
    wire __A23_1__PIPGXm;
    wire __A23_1__PIPGXp;
    wire __A23_1__PIPGYm;
    wire __A23_1__PIPGYp;
    wire __A23_1__PIPGZm;
    wire __A23_1__PIPGZp;
    wire __A23_1__PIPSAM;
    wire __A23_1__PIPSAM_n;
    wire __A23_2__CCH07;
    wire __A23_2__ISSTDC;
    wire __A23_2__OT1108;
    wire __A23_2__OT1113;
    wire __A23_2__OT1114;
    wire __A23_2__OT1116;
    wire __A23_2__RCH07_n;
    wire __A23_2__WCH07_n;
    wire __A23_NET_101;
    wire __A23_NET_102;
    wire __A23_NET_103;
    wire __A23_NET_104;
    wire __A23_NET_105;
    wire __A23_NET_106;
    wire __A23_NET_107;
    wire __A23_NET_108;
    wire __A23_NET_109;
    wire __A23_NET_110;
    wire __A23_NET_111;
    wire __A23_NET_112;
    wire __A23_NET_113;
    wire __A23_NET_114;
    wire __A23_NET_115;
    wire __A23_NET_116;
    wire __A23_NET_117;
    wire __A23_NET_118;
    wire __A23_NET_119;
    wire __A23_NET_120;
    wire __A23_NET_123;
    wire __A23_NET_126;
    wire __A23_NET_127;
    wire __A23_NET_129;
    wire __A23_NET_143;
    wire __A23_NET_144;
    wire __A23_NET_147;
    wire __A23_NET_148;
    wire __A23_NET_149;
    wire __A23_NET_153;
    wire __A23_NET_154;
    wire __A23_NET_155;
    wire __A23_NET_156;
    wire __A23_NET_157;
    wire __A23_NET_158;
    wire __A23_NET_159;
    wire __A23_NET_160;
    wire __A23_NET_161;
    wire __A23_NET_162;
    wire __A23_NET_163;
    wire __A23_NET_164;
    wire __A23_NET_165;
    wire __A23_NET_166;
    wire __A23_NET_167;
    wire __A23_NET_168;
    wire __A23_NET_169;
    wire __A23_NET_170;
    wire __A23_NET_171;
    wire __A23_NET_172;
    wire __A23_NET_173;
    wire __A23_NET_174;
    wire __A23_NET_174_U23002_6;
    wire __A23_NET_174_U23002_8;
    wire __A23_NET_175;
    wire __A23_NET_176;
    wire __A23_NET_178;
    wire __A23_NET_179;
    wire __A23_NET_182;
    wire __A23_NET_184;
    wire __A23_NET_185;
    wire __A23_NET_185_U23002_2;
    wire __A23_NET_185_U23002_4;
    wire __A23_NET_187;
    wire __A23_NET_188;
    wire __A23_NET_189;
    wire __A23_NET_190;
    wire __A23_NET_191;
    wire __A23_NET_192;
    wire __A23_NET_193;
    wire __A23_NET_194;
    wire __A23_NET_195;
    wire __A23_NET_196;
    wire __A23_NET_197;
    wire __A23_NET_198;
    wire __A23_NET_199;
    wire __A23_NET_200;
    wire __A23_NET_201;
    wire __A23_NET_202;
    wire __A23_NET_203;
    wire __A23_NET_204;
    wire __A23_NET_205;
    wire __A23_NET_206;
    wire __A23_NET_208;
    wire __A23_NET_209;
    wire __A23_NET_211;
    wire __A23_NET_212;
    wire __A23_NET_213;
    wire __A23_NET_214;
    wire __A23_NET_215;
    wire __A23_NET_216;
    wire __A23_NET_217;
    wire __A23_NET_218;
    wire __A23_NET_219;
    wire __A23_NET_220;
    wire __A23_NET_222;
    wire __A23_NET_223;
    wire __A23_NET_225;
    wire __A23_NET_227;
    wire __A23_NET_228;
    wire __A23_NET_229;
    wire __A23_NET_230;
    wire __A23_NET_231;
    wire __A23_NET_232;
    wire __A23_NET_233;
    wire __A23_NET_234;
    wire __A23_NET_235;
    wire __A23_NET_236;
    wire __A23_NET_237;
    wire __A23_NET_238;
    wire __A23_NET_239;
    wire __A23_NET_240;
    wire __A23_NET_241;
    wire __A23_NET_242;
    wire __A23_NET_243;
    wire __A23_NET_244;
    wire __A23_NET_245;
    wire __A23_NET_246;
    wire __A23_NET_247;
    wire __A23_NET_248;
    wire __A23_NET_249;
    wire __A23_NET_250;
    wire __A23_NET_251;
    wire __A23_NET_252;
    wire __A23_NET_253;
    wire __A23_NET_254;
    wire __A23_NET_255;
    wire __A23_NET_256;
    wire __A23_NET_257;
    wire __A23_NET_258;
    wire __A23_NET_259;
    wire __A23_NET_260;
    wire __A23_NET_261;
    wire __A23_NET_262;
    wire __A23_NET_263;
    wire __A23_NET_264;
    wire __A23_NET_265;
    wire __A23_NET_266;
    wire __A23_NET_267;
    wire __A23_NET_268;
    wire __A23_NET_269;
    wire __A23_NET_270;
    wire __A23_NET_271;
    wire __A23_NET_272;
    wire __A23_NET_273;
    wire __A24_1__12KPPS;
    wire __A24_1__25KPPS;
    wire __A24_1__3200A;
    wire __A24_1__3200B;
    wire __A24_1__3200C;
    wire __A24_1__3200D;
    wire __A24_1__800RST;
    wire __A24_1__800SET;
    wire __A24_1__CDUCLK;
    wire __A24_1__F03B_n;
    wire __A24_1__F07A_n;
    wire __A24_1__LRRST;
    wire __A24_1__PIPINT;
    wire __A24_1__RRRST;
    wire __A24_2__FS06_n;
    wire __A24_2__FS08_n;
    wire __A24_NET_195;
    wire __A24_NET_196;
    wire __A24_NET_197;
    wire __A24_NET_198;
    wire __A24_NET_199;
    wire __A24_NET_200;
    wire __A24_NET_201;
    wire __A24_NET_202;
    wire __A24_NET_203;
    wire __A24_NET_204;
    wire __A24_NET_205;
    wire __A24_NET_206;
    wire __A24_NET_207;
    wire __A24_NET_208;
    wire __A24_NET_209;
    wire __A24_NET_210;
    wire __A24_NET_211;
    wire __A24_NET_212;
    wire __A24_NET_213;
    wire __A24_NET_215;
    wire __A24_NET_216;
    wire __A24_NET_217;
    wire __A24_NET_219;
    wire __A24_NET_220;
    wire __A24_NET_222;
    wire __A24_NET_223;
    wire __A24_NET_226;
    wire __A24_NET_228;
    wire __A24_NET_229;
    wire __A24_NET_230;
    wire __A24_NET_233;
    wire __A24_NET_234;
    wire __A24_NET_235;
    wire __A24_NET_238;
    wire __A24_NET_239;
    wire __A24_NET_240;
    wire __A24_NET_241;
    wire __A24_NET_244;
    wire __A24_NET_245;
    wire __A24_NET_246;
    wire __A24_NET_247;
    wire __A24_NET_248;
    wire __A24_NET_249;
    wire __A24_NET_250;
    wire __A24_NET_251;
    wire __A24_NET_252;
    wire __A24_NET_253;
    wire __A24_NET_256;
    wire __B01_1__CQA;
    wire __B01_1__CQB;
    wire __B01_1__CQC;
    wire __B01_1__FADDR1;
    wire __B01_1__FADDR10;
    wire __B01_1__FADDR11;
    wire __B01_1__FADDR12;
    wire __B01_1__FADDR13;
    wire __B01_1__FADDR14;
    wire __B01_1__FADDR15;
    wire __B01_1__FADDR16;
    wire __B01_1__FADDR2;
    wire __B01_1__FADDR3;
    wire __B01_1__FADDR4;
    wire __B01_1__FADDR5;
    wire __B01_1__FADDR6;
    wire __B01_1__FADDR7;
    wire __B01_1__FADDR8;
    wire __B01_1__FADDR9;
    wire __B01_1__NOROPE;
    wire __B01_1__QUARTERA;
    wire __B01_1__QUARTERB;
    wire __B01_1__QUARTERC;
    wire __B01_2__EDESTROY;
    wire __B01_2__ES01_n;
    wire __B01_2__ES02_n;
    wire __B01_2__ES03_n;
    wire __B01_2__ES04_n;
    wire __B01_2__ES05_n;
    wire __B01_2__ES06_n;
    wire __B01_2__ES07_n;
    wire __B01_2__ES08_n;
    wire __B01_2__ES09_n;
    wire __B01_2__ES10_n;
    wire __B01_2__ES11_n;
    wire __B01_2__RADDR1;
    wire __B01_2__RADDR10;
    wire __B01_2__RADDR11;
    wire __B01_2__RADDR2;
    wire __B01_2__RADDR3;
    wire __B01_2__RADDR4;
    wire __B01_2__RADDR5;
    wire __B01_2__RADDR6;
    wire __B01_2__RADDR7;
    wire __B01_2__RADDR8;
    wire __B01_2__RADDR9;
    wire __B01_2__RESETK;
    wire __B01_NET_101;
    wire __B01_NET_103;
    wire __B01_NET_104;
    wire __B01_NET_105;
    wire __B01_NET_106;
    wire __B01_NET_107;
    wire __B01_NET_108;
    wire __B01_NET_109;
    wire __B01_NET_110;
    wire __B01_NET_111;
    wire __B01_NET_112;
    wire __B01_NET_113;
    wire __B01_NET_118;
    wire __B01_NET_123;
    wire __B01_NET_124;
    wire __B01_NET_125;
    wire __B01_NET_127;
    wire __B01_NET_128;
    wire __B01_NET_129;
    wire __B01_NET_130;
    wire __B01_NET_131;
    wire __B01_NET_133;
    wire __B01_NET_134;
    wire __B01_NET_136;
    wire __B01_NET_138;
    wire __B01_NET_139;
    wire __B01_NET_140;
    wire __B01_NET_141;
    wire __B01_NET_142;
    wire __B01_NET_143;
    wire __B01_NET_144;
    wire __B01_NET_145;
    wire __B01_NET_146;
    wire __B01_NET_147;
    wire __B01_NET_148;
    wire __B01_NET_149;
    wire __B01_NET_150;
    wire __B01_NET_152;
    wire __B01_NET_154;
    wire __B01_NET_155;
    wire __B01_NET_156;
    wire __B01_NET_157;
    wire __B01_NET_158;
    wire __B01_NET_159;
    wire __B01_NET_162;
    wire __B01_NET_166;
    wire __B01_NET_179;
    wire __B01_NET_180;
    wire __B01_NET_181;
    wire __B01_NET_184;
    wire __B01_NET_186;
    wire __B01_NET_187;
    wire __B01_NET_188;
    wire __B01_NET_189;
    wire __B01_NET_190;
    wire __B01_NET_191;
    wire __B01_NET_192;
    wire __B01_NET_194;
    wire __B01_NET_196;
    wire __B01_NET_197;
    wire __B01_NET_198;
    wire __B01_NET_199;
    wire __B01_NET_200;
    wire __B01_NET_201;
    wire __B01_NET_202;
    wire __B01_NET_203;
    wire __B01_NET_204;
    wire __B01_NET_205;
    wire __B01_NET_210;
    wire __B01_NET_211;
    wire __B01_NET_212;
    wire __B01_NET_213;
    wire __B01_NET_214;
    wire __B01_NET_215;
    wire __B01_NET_216;
    wire __B01_NET_217;
    wire __B01_NET_218;
    wire __B01_NET_220;
    wire __B01_NET_221;
    wire __B01_NET_222;
    wire __B01_NET_223;
    wire __B01_NET_224;
    wire __B01_NET_225;
    wire __B01_NET_226;
    wire __B01_NET_229;
    wire __B01_NET_230;
    wire __B01_NET_232;
    wire __B01_NET_233;
    wire __B01_NET_235;
    wire __B01_NET_236;
    wire __B01_NET_238;
    wire __B01_NET_239;
    wire __B01_NET_240;
    wire __B01_NET_241;
    wire __B01_NET_242;
    wire __B01_NET_95;
    wire __B01_NET_96;
    wire __B01_NET_98;
    wire __CG11;
    wire __CG12;
    wire __CG14;
    wire __CG21;
    wire __CG22;
    wire __CG24;
    wire __CI03_n;
    wire __CI07_n;
    wire __CI11_n;
    wire __CI15_n;
    wire __CO04;
    wire __CO04_U8007_2;
    wire __CO04_U8013_2;
    wire __CO08;
    wire __CO08_U9007_2;
    wire __CO08_U9013_2;
    wire __CO12;
    wire __CO12_U10007_2;
    wire __CO12_U10013_2;
    wire __CO16;
    wire __CO16_U11007_2;
    wire __CO16_U11013_2;
    wire __G04_n;
    wire __G04_n_U8061_10;
    wire __G04_n_U8061_12;
    wire __G08_n;
    wire __G08_n_U9061_10;
    wire __G08_n_U9061_12;
    wire __G12_n;
    wire __G12_n_U10061_10;
    wire __G12_n_U10061_12;
    wire __G16_n;
    wire __G16_n_U11061_10;
    wire __G16_n_U11061_12;
    wire __L03_n;
    wire __L03_n_U8041_6;
    wire __L05_n;
    wire __L05_n_U9007_6;
    wire __L06_n;
    wire __L06_n_U9013_12;
    wire __L07_n;
    wire __L07_n_U9041_6;
    wire __L09_n;
    wire __L09_n_U10007_6;
    wire __L10_n;
    wire __L10_n_U10013_12;
    wire __L11_n;
    wire __L11_n_U10041_6;
    wire __L13_n;
    wire __L13_n_U11007_6;
    wire __L14_n;
    wire __L14_n_U11013_12;
    wire __RL16;
    wire __XUY03_n;
    wire __XUY04_n;
    wire __XUY07_n;
    wire __XUY08_n;
    wire __XUY11_n;
    wire __XUY12_n;
    wire __XUY15_n;
    wire __XUY16_n;
    wire n10XP1;
    wire n10XP8;
    wire n11XP2;
    wire n1XP10;
    wire n2XP3;
    wire n2XP5;
    wire n2XP7;
    wire n2XP8;
    wire n3XP2;
    wire n3XP6;
    wire n3XP7;
    wire n4XP11;
    wire n4XP5;
    wire n5XP11;
    wire n5XP11_U4039_6;
    wire n5XP11_U4039_8;
    wire n5XP12;
    wire n5XP15;
    wire n5XP21;
    wire n5XP28;
    wire n5XP4;
    wire n6XP5;
    wire n6XP8;
    wire n7XP14;
    wire n7XP19;
    wire n7XP4;
    wire n7XP9;
    wire n8PP4;
    wire n8PP4_U4063_12;
    wire n8PP4_U6037_10;
    wire n8PP4_U6037_12;
    wire n8PP4_U6041_2;
    wire n8XP5;
    wire n8XP6;
    wire n9XP1;
    wire n9XP5;

    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1101(__A01_1__F02A, __A01_1__scaler_s2__FS_n, __A01_NET_176, F02B, __A01_NET_175, FS02, GND, __A01_NET_176, FS02, __A01_1__scaler_s2__FS_n, __A01_1__scaler_s2__FS_n, __A01_NET_175, FS02, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1102(__A01_1__F02A, FS01_n, __A01_NET_176, FS01_n, F02B, __A01_NET_175, GND, __A01_NET_177, __A01_1__F03A, __A01_1__F02A, __A01_NET_178, __A01_NET_176, __A01_NET_175, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1103(__A01_1__F03A, __A01_1__scaler_s3__FS_n, __A01_NET_177, F03B, __A01_NET_178, FS03, GND, __A01_NET_177, FS03, __A01_1__scaler_s3__FS_n, __A01_1__scaler_s3__FS_n, __A01_NET_178, FS03, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1104(__A01_NET_177, __A01_1__F02A, F04A, __A01_1__F03A, __A01_NET_179, __A01_NET_180, GND, __A01_NET_179, __A01_NET_180, __A01_1__F03A, F04B, __A01_NET_178, F03B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1105(F04A, __A01_1__scaler_s4__FS_n, __A01_NET_180, F04B, __A01_NET_179, FS04, GND, __A01_NET_180, FS04, __A01_1__scaler_s4__FS_n, __A01_1__scaler_s4__FS_n, __A01_NET_179, FS04, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1106(__A01_1__F05A, __A01_1__scaler_s5__FS_n, __A01_NET_181, __A01_1__F05B, __A01_NET_182, FS05, GND, __A01_NET_181, FS05, __A01_1__scaler_s5__FS_n, __A01_1__scaler_s5__FS_n, __A01_NET_182, FS05, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1107(__A01_1__F05A, F04A, __A01_NET_181, F04A, __A01_1__F05B, __A01_NET_182, GND, __A01_NET_183, __A01_1__F06A, __A01_1__F05A, __A01_NET_184, __A01_NET_181, __A01_NET_182, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1108(__A01_1__F06A, __A01_1__scaler_s6__FS_n, __A01_NET_183, F06B, __A01_NET_184, FS06, GND, __A01_NET_183, FS06, __A01_1__scaler_s6__FS_n, __A01_1__scaler_s6__FS_n, __A01_NET_184, FS06, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1109(__A01_NET_183, __A01_1__F05A, F07A, __A01_1__F06A, __A01_NET_186, __A01_NET_185, GND, __A01_NET_186, __A01_NET_185, __A01_1__F06A, F07B, __A01_NET_184, F06B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1110(F07A, __A01_1__scaler_s7__FS_n, __A01_NET_185, F07B, __A01_NET_186, __A01_1__FS07, GND, __A01_NET_185, __A01_1__FS07, __A01_1__scaler_s7__FS_n, __A01_1__scaler_s7__FS_n, __A01_NET_186, __A01_1__FS07, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1111(__A01_1__F08A, __A01_1__scaler_s8__FS_n, __A01_NET_187, F08B, __A01_NET_188, FS08, GND, __A01_NET_187, FS08, __A01_1__scaler_s8__FS_n, __A01_1__scaler_s8__FS_n, __A01_NET_188, FS08, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1112(__A01_1__F08A, F07A, __A01_NET_187, F07A, F08B, __A01_NET_188, GND, __A01_NET_189, F09A, __A01_1__F08A, __A01_NET_190, __A01_NET_187, __A01_NET_188, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1113(F09A, __A01_1__scaler_s9__FS_n, __A01_NET_189, F09B, __A01_NET_190, FS09, GND, __A01_NET_189, FS09, __A01_1__scaler_s9__FS_n, __A01_1__scaler_s9__FS_n, __A01_NET_190, FS09, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1114(__A01_NET_189, __A01_1__F08A, F10A, F09A, __A01_NET_192, __A01_NET_191, GND, __A01_NET_192, __A01_NET_191, F09A, F10B, __A01_NET_190, F09B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1115(F10A, __A01_1__scaler_s10__FS_n, __A01_NET_191, F10B, __A01_NET_192, FS10, GND, __A01_NET_191, FS10, __A01_1__scaler_s10__FS_n, __A01_1__scaler_s10__FS_n, __A01_NET_192, FS10, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1116(__A01_1__F11A, __A01_1__scaler_s11__FS_n, __A01_NET_193, __A01_1__F11B, __A01_NET_194, __A01_1__FS11, GND, __A01_NET_193, __A01_1__FS11, __A01_1__scaler_s11__FS_n, __A01_1__scaler_s11__FS_n, __A01_NET_194, __A01_1__FS11, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1117(__A01_1__F11A, F10A, __A01_NET_193, F10A, __A01_1__F11B, __A01_NET_194, GND, __A01_NET_196, __A01_1__F12A, __A01_1__F11A, __A01_NET_195, __A01_NET_193, __A01_NET_194, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1118(__A01_1__F12A, __A01_1__scaler_s12__FS_n, __A01_NET_196, F12B, __A01_NET_195, __A01_1__FS12, GND, __A01_NET_196, __A01_1__FS12, __A01_1__scaler_s12__FS_n, __A01_1__scaler_s12__FS_n, __A01_NET_195, __A01_1__FS12, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1119(__A01_NET_196, __A01_1__F11A, __A01_1__F13A, __A01_1__F12A, __A01_NET_198, __A01_NET_197, GND, __A01_NET_198, __A01_NET_197, __A01_1__F12A, __A01_1__F13B, __A01_NET_195, F12B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1120(__A01_1__F13A, __A01_1__scaler_s13__FS_n, __A01_NET_197, __A01_1__F13B, __A01_NET_198, FS13, GND, __A01_NET_197, FS13, __A01_1__scaler_s13__FS_n, __A01_1__scaler_s13__FS_n, __A01_NET_198, FS13, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1121(__A01_1__F14A, __A01_1__scaler_s14__FS_n, __A01_NET_199, F14B, __A01_NET_200, FS14, GND, __A01_NET_199, FS14, __A01_1__scaler_s14__FS_n, __A01_1__scaler_s14__FS_n, __A01_NET_200, FS14, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1122(__A01_1__F14A, __A01_1__F13A, __A01_NET_199, __A01_1__F13A, F14B, __A01_NET_200, GND, __A01_NET_202, __A01_1__F15A, __A01_1__F14A, __A01_NET_201, __A01_NET_199, __A01_NET_200, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1123(__A01_1__F15A, __A01_1__scaler_s15__FS_n, __A01_NET_202, __A01_1__F15B, __A01_NET_201, __A01_1__FS15, GND, __A01_NET_202, __A01_1__FS15, __A01_1__scaler_s15__FS_n, __A01_1__scaler_s15__FS_n, __A01_NET_201, __A01_1__FS15, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1124(__A01_NET_202, __A01_1__F14A, __A01_1__F16A, __A01_1__F15A, __A01_NET_204, __A01_NET_203, GND, __A01_NET_204, __A01_NET_203, __A01_1__F15A, __A01_1__F16B, __A01_NET_201, __A01_1__F15B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1125(__A01_1__F16A, __A01_1__scaler_s16__FS_n, __A01_NET_203, __A01_1__F16B, __A01_NET_204, FS16, GND, __A01_NET_203, FS16, __A01_1__scaler_s16__FS_n, __A01_1__scaler_s16__FS_n, __A01_NET_204, FS16, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1126(F17A, __A01_1__scaler_s17__FS_n, __A01_NET_205, F17B, __A01_NET_206, FS17, GND, __A01_NET_205, FS17, __A01_1__scaler_s17__FS_n, __A01_1__scaler_s17__FS_n, __A01_NET_206, FS17, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1127(F17A, __A01_1__F16A, __A01_NET_205, __A01_1__F16A, F17B, __A01_NET_206, GND,  ,  ,  ,  , __A01_NET_205, __A01_NET_206, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U1128(__A01_1__scaler_s2__FS_n, __A01_1__FS02A, __A01_1__scaler_s3__FS_n, __A01_1__FS03A, __A01_1__scaler_s4__FS_n, __A01_1__FS04A, GND, __A01_1__FS05A, __A01_1__scaler_s5__FS_n, F05A_n, __A01_1__F05A, F05B_n, __A01_1__F05B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1129(CHAT01, RCHAT_n, __A01_1__scaler_s6__FS_n, CHAT02, RCHAT_n, __A01_1__scaler_s7__FS_n, GND, RCHAT_n, __A01_1__scaler_s8__FS_n, CHAT03, RCHAT_n, __A01_1__scaler_s9__FS_n, CHAT04, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1130(CHAT05, RCHAT_n, __A01_1__scaler_s10__FS_n, CHAT06, RCHAT_n, __A01_1__scaler_s11__FS_n, GND, RCHAT_n, __A01_1__scaler_s12__FS_n, CHAT07, RCHAT_n, __A01_1__scaler_s13__FS_n, CHAT08, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1131(CHAT09, RCHAT_n, __A01_1__scaler_s14__FS_n, CHAT10, RCHAT_n, __A01_1__scaler_s15__FS_n, GND, RCHAT_n, __A01_1__scaler_s16__FS_n, CHAT11, RCHAT_n, __A01_1__scaler_s17__FS_n, CHAT12, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1132(F18A, __A01_2__scaler_s18__FS_n, __A01_NET_207, F18B, __A01_NET_208, __A01_2__FS18, GND, __A01_NET_207, __A01_2__FS18, __A01_2__scaler_s18__FS_n, __A01_2__scaler_s18__FS_n, __A01_NET_208, __A01_2__FS18, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1133(F18A, F17A, __A01_NET_207, F17A, F18B, __A01_NET_208, GND, __A01_NET_209, __A01_2__F19A, F18A, __A01_NET_210, __A01_NET_207, __A01_NET_208, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1134(__A01_2__F19A, __A01_2__scaler_s19__FS_n, __A01_NET_209, __A01_2__F19B, __A01_NET_210, __A01_2__FS19, GND, __A01_NET_209, __A01_2__FS19, __A01_2__scaler_s19__FS_n, __A01_2__scaler_s19__FS_n, __A01_NET_210, __A01_2__FS19, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1135(__A01_NET_209, F18A, __A01_2__F20A, __A01_2__F19A, __A01_NET_212, __A01_NET_211, GND, __A01_NET_212, __A01_NET_211, __A01_2__F19A, __A01_2__F20B, __A01_NET_210, __A01_2__F19B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1136(__A01_2__F20A, __A01_2__scaler_s20__FS_n, __A01_NET_211, __A01_2__F20B, __A01_NET_212, __A01_2__FS20, GND, __A01_NET_211, __A01_2__FS20, __A01_2__scaler_s20__FS_n, __A01_2__scaler_s20__FS_n, __A01_NET_212, __A01_2__FS20, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1137(__A01_2__F21A, __A01_2__scaler_s21__FS_n, __A01_NET_213, __A01_2__F21B, __A01_NET_214, __A01_2__FS21, GND, __A01_NET_213, __A01_2__FS21, __A01_2__scaler_s21__FS_n, __A01_2__scaler_s21__FS_n, __A01_NET_214, __A01_2__FS21, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1138(__A01_2__F21A, __A01_2__F20A, __A01_NET_213, __A01_2__F20A, __A01_2__F21B, __A01_NET_214, GND, __A01_NET_215, __A01_2__F22A, __A01_2__F21A, __A01_NET_216, __A01_NET_213, __A01_NET_214, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1139(__A01_2__F22A, __A01_2__scaler_s22__FS_n, __A01_NET_215, __A01_2__F22B, __A01_NET_216, __A01_2__FS22, GND, __A01_NET_215, __A01_2__FS22, __A01_2__scaler_s22__FS_n, __A01_2__scaler_s22__FS_n, __A01_NET_216, __A01_2__FS22, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1140(__A01_NET_215, __A01_2__F21A, __A01_2__F23A, __A01_2__F22A, __A01_NET_218, __A01_NET_217, GND, __A01_NET_218, __A01_NET_217, __A01_2__F22A, __A01_2__F23B, __A01_NET_216, __A01_2__F22B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1141(__A01_2__F23A, __A01_2__scaler_s23__FS_n, __A01_NET_217, __A01_2__F23B, __A01_NET_218, __A01_2__FS23, GND, __A01_NET_217, __A01_2__FS23, __A01_2__scaler_s23__FS_n, __A01_2__scaler_s23__FS_n, __A01_NET_218, __A01_2__FS23, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1142(__A01_2__F24A, __A01_2__scaler_s24__FS_n, __A01_NET_219, __A01_2__F24B, __A01_NET_220, __A01_2__FS24, GND, __A01_NET_219, __A01_2__FS24, __A01_2__scaler_s24__FS_n, __A01_2__scaler_s24__FS_n, __A01_NET_220, __A01_2__FS24, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1143(__A01_2__F24A, __A01_2__F23A, __A01_NET_219, __A01_2__F23A, __A01_2__F24B, __A01_NET_220, GND, __A01_NET_221, __A01_2__F25A, __A01_2__F24A, __A01_NET_222, __A01_NET_219, __A01_NET_220, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1144(__A01_2__F25A, __A01_2__scaler_s25__FS_n, __A01_NET_221, __A01_2__F25B, __A01_NET_222, __A01_2__FS25, GND, __A01_NET_221, __A01_2__FS25, __A01_2__scaler_s25__FS_n, __A01_2__scaler_s25__FS_n, __A01_NET_222, __A01_2__FS25, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1145(__A01_NET_221, __A01_2__F24A, __A01_2__F26A, __A01_2__F25A, __A01_NET_224, __A01_NET_223, GND, __A01_NET_224, __A01_NET_223, __A01_2__F25A, __A01_2__F26B, __A01_NET_222, __A01_2__F25B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1146(__A01_2__F26A, __A01_2__scaler_s26__FS_n, __A01_NET_223, __A01_2__F26B, __A01_NET_224, __A01_2__FS26, GND, __A01_NET_223, __A01_2__FS26, __A01_2__scaler_s26__FS_n, __A01_2__scaler_s26__FS_n, __A01_NET_224, __A01_2__FS26, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1147(__A01_2__F27A, __A01_2__scaler_s27__FS_n, __A01_NET_225, __A01_2__F27B, __A01_NET_226, __A01_2__FS27, GND, __A01_NET_225, __A01_2__FS27, __A01_2__scaler_s27__FS_n, __A01_2__scaler_s27__FS_n, __A01_NET_226, __A01_2__FS27, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1148(__A01_2__F27A, __A01_2__F26A, __A01_NET_225, __A01_2__F26A, __A01_2__F27B, __A01_NET_226, GND, __A01_NET_227, __A01_2__F28A, __A01_2__F27A, __A01_NET_228, __A01_NET_225, __A01_NET_226, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1149(__A01_2__F28A, __A01_2__scaler_s28__FS_n, __A01_NET_227, __A01_2__F28B, __A01_NET_228, __A01_2__FS28, GND, __A01_NET_227, __A01_2__FS28, __A01_2__scaler_s28__FS_n, __A01_2__scaler_s28__FS_n, __A01_NET_228, __A01_2__FS28, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1150(__A01_NET_227, __A01_2__F27A, __A01_2__F29A, __A01_2__F28A, __A01_NET_230, __A01_NET_229, GND, __A01_NET_230, __A01_NET_229, __A01_2__F28A, __A01_2__F29B, __A01_NET_228, __A01_2__F28B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1151(__A01_2__F29A, __A01_2__scaler_s29__FS_n, __A01_NET_229, __A01_2__F29B, __A01_NET_230, __A01_2__FS29, GND, __A01_NET_229, __A01_2__FS29, __A01_2__scaler_s29__FS_n, __A01_2__scaler_s29__FS_n, __A01_NET_230, __A01_2__FS29, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1152(__A01_2__F30A, __A01_2__scaler_s30__FS_n, __A01_NET_231, __A01_2__F30B, __A01_NET_232, __A01_2__FS30, GND, __A01_NET_231, __A01_2__FS30, __A01_2__scaler_s30__FS_n, __A01_2__scaler_s30__FS_n, __A01_NET_232, __A01_2__FS30, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1153(__A01_2__F30A, __A01_2__F29A, __A01_NET_231, __A01_2__F29A, __A01_2__F30B, __A01_NET_232, GND, __A01_NET_233, __A01_2__F31A, __A01_2__F30A, __A01_NET_234, __A01_NET_231, __A01_NET_232, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1154(__A01_2__F31A, __A01_2__scaler_s31__FS_n, __A01_NET_233, __A01_2__F31B, __A01_NET_234, __A01_2__FS31, GND, __A01_NET_233, __A01_2__FS31, __A01_2__scaler_s31__FS_n, __A01_2__scaler_s31__FS_n, __A01_NET_234, __A01_2__FS31, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1155(__A01_NET_233, __A01_2__F30A, __A01_2__F32A, __A01_2__F31A, __A01_NET_236, __A01_NET_235, GND, __A01_NET_236, __A01_NET_235, __A01_2__F31A, __A01_2__F32B, __A01_NET_234, __A01_2__F31B, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1156(__A01_2__F32A, __A01_2__scaler_s32__FS_n, __A01_NET_235, __A01_2__F32B, __A01_NET_236, __A01_2__FS32, GND, __A01_NET_235, __A01_2__FS32, __A01_2__scaler_s32__FS_n, __A01_2__scaler_s32__FS_n, __A01_NET_236, __A01_2__FS32, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U1157(__A01_2__F33A, __A01_2__scaler_s33__FS_n, __A01_NET_237, __A01_2__F33B, __A01_NET_238, __A01_2__FS33, GND, __A01_NET_237, __A01_2__FS33, __A01_2__scaler_s33__FS_n, __A01_2__scaler_s33__FS_n, __A01_NET_238, __A01_2__FS33, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U1158(__A01_2__F33A, __A01_2__F32A, __A01_NET_237, __A01_2__F32A, __A01_2__F33B, __A01_NET_238, GND,  ,  ,  ,  , __A01_NET_237, __A01_NET_238, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1159(CHAT13, RCHAT_n, __A01_2__scaler_s18__FS_n, CHAT14, RCHAT_n, __A01_2__scaler_s19__FS_n, GND, RCHBT_n, __A01_2__scaler_s20__FS_n, CHBT01, RCHBT_n, __A01_2__scaler_s21__FS_n, CHBT02, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1160(CHBT03, RCHBT_n, __A01_2__scaler_s22__FS_n, CHBT04, RCHBT_n, __A01_2__scaler_s23__FS_n, GND, RCHBT_n, __A01_2__scaler_s24__FS_n, CHBT05, RCHBT_n, __A01_2__scaler_s25__FS_n, CHBT06, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1161(CHBT07, RCHBT_n, __A01_2__scaler_s26__FS_n, CHBT08, RCHBT_n, __A01_2__scaler_s27__FS_n, GND, RCHBT_n, __A01_2__scaler_s28__FS_n, CHBT09, RCHBT_n, __A01_2__scaler_s29__FS_n, CHBT10, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U1162(CHBT11, RCHBT_n, __A01_2__scaler_s30__FS_n, CHBT12, RCHBT_n, __A01_2__scaler_s31__FS_n, GND, RCHBT_n, __A01_2__scaler_s32__FS_n, CHBT13, RCHBT_n, __A01_2__scaler_s33__FS_n, CHBT14, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U1163(F07B, F07B_n, F10A, F10A_n, F09B, F09B_n, GND, FS07_n, __A01_1__FS07, FS07A, FS07_n, FS05_n, FS05, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U1164(FS09, FS09_n,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2101(__A02_1__cdiv_1__D, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__B, __A02_1__cdiv_1__FS, GND, __A02_1__cdiv_1__FS_n, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, __A02_1__cdiv_1__A, __A02_1__cdiv_1__FS, PHS2, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U2102(__A02_1__cdiv_1__D, CLOCK, __A02_1__cdiv_1__B, CLOCK, PHS2, __A02_1__cdiv_1__A, GND, __A02_2__EDSET, P02, P03_n, P04, __A02_1__cdiv_1__B, __A02_1__cdiv_1__A, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1) U2103(__A02_1__cdiv_1__D, __A02_1__cdiv_2__F, PHS2, PHS2_n, PHS4, PHS4_n, GND, __A02_NET_133, __A02_1__cdiv_1__B, CT, __A02_NET_133, CT_n, CT, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U2104(PHS4, __A02_1__cdiv_2__F, __A02_1__cdiv_1__A, __A02_1__oddset, STOP, __A02_1__RINGA_n, GND, P02_n, P04, SB4, P02_n, P05, __A02_2__SB0, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1) U2105(__A02_1__cdiv_1__FS_n, WT, WT, WT_n, WT, TT_n, GND, __A02_1__ovfstb_r5, __A02_1__ovfstb_r4, __A02_1__ovfstb_r6, __A02_1__ovfstb_r5, __A02_1__OVFSTB_n, __A02_1__ovfstb_r2, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2106(__A02_1__cdiv_2__D, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__FS, GND, __A02_1__cdiv_2__FS_n, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__A, __A02_1__cdiv_2__FS, __A02_1__cdiv_2__C, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U2107(__A02_1__cdiv_2__D, __A02_1__cdiv_2__F, __A02_1__cdiv_2__B, __A02_1__cdiv_2__F, __A02_1__cdiv_2__C, __A02_1__cdiv_2__A, GND, P03, __A02_2__EDSET, __A02_NET_158, P03_n, __A02_1__cdiv_2__B, __A02_1__cdiv_2__A, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U2108(__A02_1__cdiv_2__D, __A02_1__RINGA_n, __A02_1__oddset, __A02_1__ODDSET_n, __A02_1__cdiv_2__C, __A02_1__RINGB_n, GND, __A02_1__evnset, __A02_1__RINGB_n, __A02_1__EVNSET_n, __A02_1__evnset, RT, __A02_1__cdiv_1__A, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U2109(__A02_1__ovfstb_r1, CT_n, __A02_1__ovfstb_r2, __A02_1__ovfstb_r2, __A02_1__ovfstb_r6, __A02_1__ovfstb_r1, GND, __A02_1__ovfstb_r4, __A02_1__ovfstb_r2, __A02_1__ovfstb_r3, __A02_1__ovfstb_r3, __A02_1__ovfstb_r1, __A02_1__ovfstb_r4, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U2110(CT, PHS3_n, WT_n, CLK,  ,  , GND,  ,  , RT_n, RT,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U2111(__A02_1__RINGB_n, P05_n, P04, P05, __A02_1__RINGA_n, __A02_NET_162, GND, __A02_NET_143, __A02_2__T12DC_n, __A02_NET_151, __A02_1__EVNSET_n, __A02_NET_163, P04_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2112(P01, __A02_NET_163, P01_n, P01_n, P01, __A02_NET_162, GND, __A02_1__RINGA_n, P01, __A02_NET_168, P01_n, __A02_1__RINGB_n, __A02_NET_167, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2113(P02, __A02_NET_168, P02_n, P02_n, P02, __A02_NET_167, GND, __A02_1__RINGB_n, P02, __A02_NET_158, P02_n, __A02_1__RINGA_n, __A02_NET_166, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2114(__A02_2__SB1, P05_n, P03_n, P03_n, P03, __A02_NET_166, GND, __A02_1__RINGA_n, P03, __A02_NET_170, P03_n, __A02_1__RINGB_n, __A02_NET_169, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2115(P04, __A02_NET_170, P04_n, P04_n, P04, __A02_NET_169, GND, __A02_1__RINGB_n, P04, __A02_NET_165, P04_n, __A02_1__RINGA_n, __A02_NET_164, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2116(P05, __A02_NET_165, P05_n, P05_n, P05, __A02_NET_164, GND, __A02_NET_151, GOJ1, __A02_NET_154, __A02_1__EVNSET_n, __A02_NET_149, __A02_NET_144, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2117(__A02_2__F01D, FS01_n, F01B, FS01_n, F01B, FS01, GND, FS01_n, F01A, FS01, F01A, FS01, __A02_2__F01C, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U2118(__A02_2__F01D, P01_n, F01B, P01_n, __A02_2__F01C, F01A, GND,  ,  ,  ,  , F01B, F01A, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b1, 1'b0) U2119(SBY, ALGA, STRT1, STRT2, __A02_NET_154, __A02_NET_152, GND, __A02_NET_148, __A02_2__T12DC_n, __A02_NET_153, __A02_1__EVNSET_n, __A02_NET_150, MSTRTP, p4VDC, SIM_RST, SIM_CLK);
    U74LVC07 U2120(__A02_NET_150, __A02_NET_151_U2120_2, __A02_NET_152, __A02_NET_151_U2120_4,  ,  , GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0) U2121(__A02_NET_151, __A02_NET_149, MSTP, __A02_NET_153, GOJAM_n, GOJAM, GND,  ,  , STOP, STOP_n,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U2122(__A02_NET_146, __A02_1__EVNSET_n, MSTP, GOJAM_n, STRT2, STOPA, GND, STOPA, __A02_NET_145, STOP_n, P05_n, P02, SB2, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U2123(__A02_NET_142, __A02_NET_143, STOPA, STOPA, __A02_NET_142, __A02_NET_144, GND, __A02_NET_148, __A02_NET_145, __A02_NET_147, __A02_NET_147, __A02_NET_146, __A02_NET_145, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U2024(__A02_3__T12SET, GOJAM, __A02_3__T01DC_n, __A02_NET_192, GOJAM, __A02_NET_191, GND, __A02_NET_192, __A02_3__T02DC_n, __A02_NET_193, GOJAM, __A02_2__T12DC_n, __A02_NET_194, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U2025(__A02_NET_194, __A02_2__T12DC_n, __A02_NET_191, __A02_NET_195, __A02_2__T12DC_n, __A02_1__ODDSET_n, GND, __A02_2__T12DC_n, __A02_1__EVNSET_n, T12, __A02_NET_195, __A02_NET_191, __A02_3__T01DC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U2026(__A02_NET_198, __A02_3__T01DC_n, __A02_1__EVNSET_n, T01, __A02_3__T01DC_n, __A02_1__ODDSET_n, GND, __A02_NET_198, __A02_NET_192, __A02_3__T02DC_n, __A02_3__T02DC_n, __A02_1__ODDSET_n, __A02_NET_179, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2027(T02, __A02_3__T02DC_n, __A02_1__EVNSET_n, __A02_3__T03DC_n, __A02_NET_179, __A02_NET_193, GND, __A02_3__T03DC_n, __A02_1__EVNSET_n, __A02_NET_180, __A02_3__T03DC_n, __A02_1__ODDSET_n, T03, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U2028(__A02_3__T03DC_n, __A02_NET_196, __A02_3__T04DC_n, __A02_NET_197, GOJAM, __A02_NET_196, GND, __A02_NET_197, __A02_3__T05DC_n, __A02_NET_188, GOJAM, __A02_NET_193, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U2029(__A02_3__T04DC_n, __A02_NET_180, __A02_NET_196, __A02_NET_177, __A02_3__T04DC_n, __A02_1__ODDSET_n, GND, __A02_3__T04DC_n, __A02_1__EVNSET_n, T04, __A02_NET_177, __A02_NET_197, __A02_3__T05DC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U2030(__A02_NET_171, __A02_3__T05DC_n, __A02_1__EVNSET_n, T05, __A02_3__T05DC_n, __A02_1__ODDSET_n, GND, __A02_NET_188, __A02_NET_171, __A02_3__T06DC_n, __A02_1__EVNSET_n, __A02_3__T06DC_n, T06, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U2031(GOJAM, __A02_NET_186, GOJAM, __A02_NET_187, __A02_3__T07DC_n, __A02_NET_186, GND, __A02_NET_187, GOJAM, __A02_NET_190, __A02_3__T08DC_n, __A02_NET_188, __A02_3__T06DC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2032(__A02_NET_178, __A02_1__ODDSET_n, __A02_3__T06DC_n, __A02_3__T07DC_n, __A02_NET_186, __A02_NET_178, GND, __A02_1__ODDSET_n, __A02_3__T07DC_n, T07, __A02_1__EVNSET_n, __A02_3__T07DC_n, __A02_NET_184, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U2033(__A02_3__T08DC_n, __A02_NET_187, __A02_NET_184, T08, __A02_1__EVNSET_n, __A02_3__T08DC_n, GND, __A02_1__ODDSET_n, __A02_3__T08DC_n, __A02_NET_185, __A02_NET_190, __A02_NET_185, __A02_3__T09DC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U2034(GOJAM, __A02_NET_189, GOJAM, __A02_NET_199, __A02_3__T10DC_n, __A02_NET_189, GND, __A02_NET_199, GOJAM, __A02_NET_183, __A02_NET_176, __A02_NET_190, __A02_3__T09DC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U2035(T09, __A02_1__ODDSET_n, __A02_3__T09DC_n, __A02_NET_182, __A02_1__EVNSET_n, __A02_3__T09DC_n, GND, __A02_NET_189, __A02_NET_182, __A02_3__T10DC_n, __A02_1__EVNSET_n, __A02_NET_189, __A02_NET_183, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U2036(__A02_NET_181, __A02_1__ODDSET_n, __A02_3__T10DC_n, __A02_NET_176, __A02_NET_199, __A02_NET_181, GND, __A02_1__EVNSET_n, __A02_3__T10DC_n, T10, __A02_1__ODDSET_n, __A02_NET_176, T11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U2037(__A02_NET_197, __A02_NET_196, __A02_NET_190, __A02_NET_189, __A02_1__EVNSET_n, __A02_NET_174, GND, __A02_NET_175, __A02_NET_188, __A02_NET_186, __A02_NET_187, __A02_NET_173, __A02_NET_193, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U2038(__A02_NET_172, __A02_3__T12SET_U2038_2, __A02_NET_173, __A02_3__T12SET_U2038_4, __A02_NET_174, __A02_3__T12SET_U2038_6, GND, __A02_3__T12SET_U2038_8, __A02_NET_175,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1) U2039(T01, T01_n, T02, T02_n, T03, T03_n, GND, T04_n, T04, T05_n, T05, T06_n, T06, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1) U2040(T07, T07_n, T08, T08_n, T09, T09_n, GND, T10_n, T10, T11_n, T11, T12_n, T12, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U2041(WL15_n, WL16, __A02_1__OVFSTB_n, WL15, WL16_n, __A02_3__UNF, GND,  ,  ,  ,  , __A02_3__OVF, __A02_1__OVFSTB_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U2042(__A02_3__OVF, OVF_n, __A02_3__UNF, UNF_n, T12_n, T12A, GND, TIMR, __A02_NET_160,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U2043(__A02_NET_161, P04, P05_n, __A02_NET_156, STOP_n,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U2044(__A02_NET_172, __A02_NET_192, __A02_NET_191, __A02_NET_156, P01, __A02_NET_159, GND, __A02_NET_156, STOP_n, __A02_NET_159, STRT2, __A02_NET_161, __A02_NET_160, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0) U2145(__A02_2__SB0, SB0_n, __A02_2__SB1, SB1_n, SB2, SB2_n, GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74LVC06 U2046(T01_n, MT01_U2046_2, T02_n, MT02_U2046_4, T03_n, MT03_U2046_6, GND, MT04_U2046_8, T04_n, MT05_U2046_10, T05_n, MT06_U2046_12, T06_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U2047(T07_n, MT07_U2047_2, T08_n, MT08_U2047_4, T09_n, MT09_U2047_6, GND, MT10_U2047_8, T10_n, MT11_U2047_10, T11_n, MT12_U2047_12, T12_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U2148(WT_n, MONWT_U2148_2, WT_n, __A02_1__Q2A_U2148_4, GOJAM_n, MGOJAM_U2148_6, GND, MSTPIT_n_U2148_8, STOP,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U3001(__A03_NET_211, NISQ, __A03_1__NISQL, __A03_NET_213, STRTFC, __A03_NET_220, GND, RT_n, __A03_NET_209, RBSQ, __A03_NET_209, WT_n, __A03_1__wsqg, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3002(__A03_NET_211, __A03_1__INKBT1, T12_n, __A03_NET_211, __A03_1__RPTFRC, __A03_NET_220, GND, __A03_1__CSQG, T12_n, CT_n, __A03_NET_213, __A03_1__NISQL, STRTFC, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1) U3003(__A03_1__NISQL, NISQL_n, __A03_NET_220, __A03_NET_209, __A03_1__wsqg, __A03_1__WSQG_n, GND, STRTFC, __A03_NET_217, SQEXT, __A03_NET_216, SQEXT_n, __A03_NET_221, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U3004(__A03_NET_165, WL16_n, __A03_1__WSQG_n, __A03_NET_166, WL14_n, __A03_1__WSQG_n, GND, WL13_n, __A03_1__WSQG_n, __A03_NET_167, __A03_NET_190, __A03_NET_187, __A03_NET_185, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3005(__A03_NET_217, GOJAM, MTCSAI, __A03_NET_218, NISQL_n, T12_n, GND, STRTFC, __A03_NET_218, __A03_NET_219, __A03_NET_219, __A03_NET_182, __A03_NET_215, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U3006(EXTPLS, EXT, __A03_NET_182, __A03_1__INKBT1, STRTFC, FUTEXT, GND, __A03_NET_216, __A03_1__RPTFRC, __A03_NET_215, __A03_NET_221, __A03_NET_182, FUTEXT, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U3007(__A03_NET_214, __A03_NET_219, FUTEXT, __A03_NET_221, __A03_NET_216, __A03_NET_214, GND, INHPLS, __A03_1__INHINT, __A03_NET_180, KRPT, IIP, IIP_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3009(__A03_NET_180, RELPLS, IIP_n, GOJAM, n5XP4, IIP, GND, __A03_NET_178, FUTEXT, NISQL_n, T12_n, __A03_1__INHINT, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3010(PHS2_n, RUPTOR_n, __A03_1__OVNHRP, __A03_1__INHINT, IIP, __A03_NET_177, GND, __A03_NET_183, __A03_NET_181, STRTFC, T02, __A03_NET_179, MNHRPT, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U3011(__A03_NET_178, RPTSET_U3011_2, __A03_NET_179, RPTSET_U3011_4, __A03_NET_177, RPTSET_U3011_6, GND, __A03_2__IC13_n_U3011_8, __A03_NET_238, __A03_2__IC13_n_U3011_10, __A03_NET_239,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b1) U3012(__A03_NET_181, RPTSET, __A03_NET_183, __A03_NET_192, __A03_NET_165, __A03_1__SQR16, GND, __A03_NET_166, __A03_1__SQR14, __A03_NET_193, __A03_NET_167, __A03_1__SQR13, __A03_NET_194, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3013(__A03_NET_192, __A03_1__RPTFRC, __A03_NET_193, __A03_1__RPTFRC, __A03_1__CSQG, __A03_1__SQR14, GND, __A03_1__SQR13, __A03_NET_194, __A03_1__RPTFRC, __A03_1__CSQG, __A03_1__SQR16, __A03_1__CSQG, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U3014(__A03_NET_163, __A03_NET_192, INKL, __A03_NET_164, INKL, __A03_1__SQR16, GND, __A03_NET_184, __A03_1__OVNHRP, __A03_NET_189, __A03_NET_185, NISQ_n, __A03_NET_184, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U3015(__A03_NET_198, __A03_NET_168, __A03_NET_194, __A03_NET_168, __A03_NET_175, __A03_NET_169, GND, __A03_NET_170, __A03_NET_198, __A03_NET_193, __A03_NET_175, __A03_NET_176, __A03_NET_175, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3016(__A03_NET_194, __A03_NET_193, __A03_NET_198, __A03_NET_168, __A03_NET_199, __A03_NET_172, GND, __A03_NET_204, __A03_NET_194, __A03_NET_168, __A03_NET_199, __A03_NET_171, __A03_NET_175, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U3017(__A03_NET_198, __A03_NET_199, __A03_NET_194, __A03_NET_193, __A03_NET_199, __A03_NET_174, GND, __A03_NET_205, __A03_1__RPTFRC, __A03_NET_200, __A03_1__SQR12, __A03_NET_173, __A03_NET_193, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3018(__A03_NET_169, SQ1_n, __A03_NET_170, SQ2_n, __A03_NET_171, __A03_1__SQ3_n, GND, __A03_1__SQ4_n, __A03_NET_172, __A03_1__SQ6_n, __A03_NET_173, __A03_1__SQ7_n, __A03_NET_174, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3019(__A03_NET_200, WL12_n, __A03_1__WSQG_n, __A03_NET_197, WL11_n, __A03_1__WSQG_n, GND, __A03_NET_205, __A03_1__CSQG, __A03_1__SQR12, __A03_NET_196, __A03_1__CSQG, __A03_1__SQR11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b1, 1'b0) U3020(__A03_1__RPTFRC, __A03_NET_197, __A03_1__RPTFRC, __A03_NET_201, __A03_NET_202, __A03_NET_203, GND, __A03_1__INKBT1, INKL, T01_n, STD2, __A03_NET_196, __A03_1__SQR11, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3021(A16_n, __A03_NET_188, A15_n, __A03_NET_186,  ,  , GND, SQR12_n, __A03_1__SQR12, __A03_1__RPTFRC, __A03_NET_181, __A03_1__SQ5_n, __A03_NET_204, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3022(__A03_1__QC0, __A03_1__SQR11, __A03_1__SQR12, __A03_NET_206, __A03_NET_196, __A03_1__SQR12, GND, __A03_1__SQR11, __A03_NET_205, __A03_NET_207, __A03_NET_205, __A03_NET_196, __A03_NET_208, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3023(__A03_1__QC0, QC0_n, __A03_NET_206, QC1_n, __A03_NET_207, QC2_n, GND, QC3_n, __A03_NET_208, SQR10, __A03_NET_203, SQR10_n, __A03_NET_202, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3024(__A03_NET_201, WL10_n, __A03_1__WSQG_n, __A03_NET_202, __A03_NET_203, __A03_1__CSQG, GND, __A03_NET_188, A15_n, __A03_NET_190, A16_n, __A03_NET_186, __A03_NET_187, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3025(__A03_NET_163, __A03_NET_199, __A03_NET_164, __A03_NET_175, __A03_NET_193, __A03_NET_168, GND, __A03_NET_198, __A03_NET_194, SQ0_n, __A03_NET_176, MP3A, MP3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3026(__A03_NET_235, __A03_1__SQ5_n, QC0_n, __A03_NET_236, __A03_1__SQ5_n, SQEXT_n, GND, __A03_NET_235, __A03_NET_236, __A03_NET_242, __A03_NET_242, ST0_n, IC1, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1) U3027(__A03_NET_235, __A03_2__SQ5QC0_n, IC2, IC2_n, __A03_NET_228, EXST1_n, GND, TC0_n, TC0, IC3, __A03_2__IC3_n, __A03_2__NEXST0_n, __A03_2__NEXST0, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3028(IC2, __A03_NET_242, ST1_n, __A03_NET_237, SQEXT_n, __A03_1__QC0, GND, SQEXT_n, ST1_n, __A03_NET_228, __A03_NET_228, __A03_2__NEXST0, __A03_NET_234, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3029(__A03_NET_237, __A03_1__SQ6_n, SQ1_n, __A03_2__NEXST0_n, __A03_1__QC0, TCF0, GND, __A03_2__IC3_n, TC0, STD2, TCF0, IC11, ST0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3030(IC6, __A03_NET_234, __A03_1__SQ3_n, IC7, __A03_NET_234, __A03_1__SQ4_n, GND, SQ0_n, __A03_2__NEXST0_n, TC0, SQEXT, ST0_n, __A03_2__NEXST0, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3031(DCS0, __A03_1__SQ4_n, EXST0_n, DCA0, EXST0_n, __A03_1__SQ3_n, GND, DCS0, DCA0, __A03_2__IC4_n, QC1_n, ST1_n, __A03_NET_240, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3032(IC7, IC6, IC1, DCS0, DCA0, __A03_NET_239, GND, IC5, __A03_NET_231, __A03_1__SQ5_n, SQEXT, __A03_NET_238, IC11, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3033(__A03_2__IC4_n, IC4, __A03_2__IC13_n, IC13, IC5, IC5_n, GND, IC9, __A03_2__IC9_n, QXCH0_n, __A03_2__QXCH0, EXST0_n, __A03_NET_223, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3034(__A03_NET_232, QC3_n, ST0_n, __A03_NET_231, __A03_NET_240, __A03_NET_232, GND, __A03_2__LXCH0, DXCH0, IC8_n, ST0_n, SQEXT_n, __A03_NET_223, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3035(__A03_2__NEXST0_n, QC1_n, SQ2_n, QC1_n, EXST0_n, __A03_2__QXCH0, GND, TS0, __A03_1__SQ5_n, QC2_n, __A03_2__NEXST0_n, __A03_2__LXCH0, SQ2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U3036(__A03_2__IC9_n, IC5, TS0, __A03_2__QXCH0, __A03_2__LXCH0,  , GND,  , SQ2_n, QC0_n, SQEXT, ST1_n, __A03_NET_224, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3037(TS0, TS0_n, IC10_n, IC10, DAS0, DAS0_n, GND, __A03_2__BZF0_n, __A03_2__BZF0, __A03_2__BMF0_n, __A03_2__BMF0, IC16, IC16_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3038(__A03_1__SQ5_n, __A03_2__NEXST0_n, SQ2_n, __A03_2__NEXST0_n, QC0_n, DAS0, GND, IC10_n, IC4, DXCH0, DAS0, DXCH0, QC1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3039(SQ1_n, __A03_1__QC0, EXST0_n, __A03_1__QC0, __A03_1__SQ6_n, __A03_2__BMF0, GND, CCS0, SQ1_n, QC0_n, __A03_2__NEXST0_n, __A03_2__BZF0, EXST0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3040(IC15_n, __A03_2__BMF0, __A03_2__BZF0, __A03_NET_226, __A03_2__BZF0_n, BR2_n, GND, __A03_2__BMF0_n, BR1B2B, __A03_NET_225, __A03_NET_226, __A03_NET_225, IC16_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U3041(IC17, IC16, IC15_n, DAS1_n, __A03_NET_224, ADS0, GND, CCS0, MSU0, IC12_n, __A03_1__SQ7_n, __A03_2__NEXST0_n, MASK0, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3042(IC15_n, IC15, CCS0, CCS0_n, DAS1_n, DAS1, GND, IC12, IC12_n, MSU0_n, MSU0, AUG0_n, __A03_2__AUG0, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U3043(SQ2_n, QC3_n, QC2_n, SQ2_n, __A03_2__NEXST0_n, INCR0, GND, MSU0, SQ2_n, EXST0_n, QC0_n, ADS0, __A03_2__NEXST0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3044(SQ2_n, EXST0_n, SQ2_n, EXST0_n, QC3_n, __A03_2__DIM0, GND, MP3, ST3_n, __A03_1__SQ7_n, SQEXT_n, __A03_2__AUG0, QC2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U3045(__A03_2__DIM0, DIM0_n, MP3, MP3_n, MP1, MP1_n, GND, MP0_n, MP0, TCSAJ3_n, TCSAJ3, RSM3_n, RSM3, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3046(ST1_n, __A03_1__SQ7_n, ST0_n, __A03_1__SQ7_n, SQEXT_n, MP0, GND, TCSAJ3, SQ0_n, SQEXT, ST3_n, MP1, SQEXT_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3047(ST3_n, __A03_2__SQ5QC0_n, __A03_1__SQ6_n, EXST0_n, QC0_n, SU0, GND, __A03_NET_227, MP0, MASK0, RXOR0, RSM3, SQEXT, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U3048(MASK0, MASK0_n, __A03_NET_227, IC14, __A03_2__NDX0, NDX0_n, GND, NDXX1_n, __A03_2__NDXX1, GOJ1_n, GOJ1, IC11_n, IC11, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U3049(AD0, __A03_2__NEXST0_n, __A03_1__SQ6_n,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3050(__A03_2__NEXST0_n, __A03_1__SQ5_n, SQEXT_n, __A03_1__SQ5_n, ST1_n, __A03_2__NDXX1, GND, GOJ1, SQEXT, ST1_n, SQ0_n, __A03_2__NDX0, QC0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U3052(__A03_NET_189, __A03_NET_191, __A03_NET_190, __A03_NET_187, NISQ_n, __A03_NET_191, GND,  ,  ,  ,  , __A03_1__OVNHRP, MP3, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U3053(__A03_NET_203, MSQ10_U3053_2, __A03_NET_180, MINHL_U3053_4, IIP_n, MIIP_U3053_6, GND, MTCSA_n_U3053_8, TCSAJ3,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U3054(__A03_NET_216, MSQEXT_U3054_2, __A03_NET_192, MSQ16_U3054_4, __A03_NET_193, MSQ14_U3054_6, GND, MSQ13_U3054_8, __A03_NET_194, MSQ12_U3054_10, __A03_NET_205, MSQ11_U3054_12, __A03_NET_196, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U4001(T12USE_n, DVST, __A04_NET_245, DIVSTG, T12USE_n, T03_n, GND, __A04_NET_247, __A04_NET_246, __A04_NET_261, GOJAM, MTCSAI, __A04_NET_252, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U4002(T03_n, T12USE_n, T12USE_n, RSTSTG, GOJAM, __A04_NET_245, GND, __A04_NET_246, PHS3_n, __A04_NET_245, T12_n, __A04_NET_247, PHS3_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U4003(__A04_NET_252, __A04_NET_249_U4003_2, __A04_NET_253, __A04_NET_249_U4003_4, __A04_NET_234, __A04_NET_236_U4003_6, GND, __A04_NET_236_U4003_8, __A04_NET_232, __A04_1__SGUM_U4003_10, __A04_NET_200, __A04_1__SGUM_U4003_12, __A04_NET_201, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b1, 1'b0) U4004(ST1, __A04_NET_248, __A04_1__STG1, __A04_1__STG3, __A04_1__STG2, __A04_NET_235, GND, __A04_NET_256, __A04_1__STG2, __A04_1__STG3, __A04_NET_244, __A04_NET_253, __A04_NET_237, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4005(__A04_NET_237, __A04_NET_249, T01, __A04_NET_248, __A04_1__DVST_n, __A04_1__STG3, GND, __A04_NET_261, __A04_NET_249, __A04_NET_250, __A04_NET_237, __A04_NET_261, __A04_NET_251, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U4006(__A04_NET_244, __A04_NET_250, __A04_1__STG1, __A04_1__STG1, __A04_NET_244, __A04_NET_251, GND, ST2, __A04_NET_241, __A04_NET_234, __A04_1__DVST_n, __A04_NET_244, __A04_NET_231, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0) U4008(__A04_NET_235, ST0_n, __A04_NET_256, ST1_n, __A04_NET_266, ST3_n, GND, __A04_1__ST4_n, __A04_NET_258, __A04_1__ST376_n, __A04_1__ST376, DV1376_n, DV1376, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U4009(__A04_NET_231, MTCSAI, __A04_NET_236, GOJAM, T01, __A04_NET_233, GND, __A04_NET_266, __A04_1__STG3, __A04_NET_257, __A04_NET_244, __A04_NET_232, __A04_NET_233, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U4010(__A04_NET_241, __A04_1__TRSM_n, XT1_n, XB7_n, NDR100_n,  , GND,  , __A04_NET_262, STRTFC, T01, RSTSTG, __A04_NET_263, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U4011(__A04_NET_238, __A04_NET_261, __A04_NET_236, __A04_NET_239, __A04_NET_233, __A04_NET_261, GND, __A04_NET_238, __A04_1__STG2, __A04_NET_257, __A04_NET_257, __A04_NET_239, __A04_1__STG2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U4012(__A04_NET_260, __A04_1__DVST_n, __A04_NET_257, __A04_NET_262, __A04_NET_260, __A04_NET_263, GND, __A04_NET_261, __A04_NET_262, __A04_NET_269, __A04_NET_263, __A04_NET_261, __A04_NET_270, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U4013(__A04_NET_214, __A04_NET_269, __A04_1__STG3, __A04_1__STG3, __A04_NET_214, __A04_NET_270, GND, __A04_1__STG1, __A04_1__STG3, __A04_NET_254, __A04_NET_257, __A04_NET_254, __A04_1__ST376, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U4014(STD2, INKL, __A04_1__STG1, __A04_1__STG3, __A04_NET_257,  , GND,  , SQ0_n, EXST1_n, QC3_n, SQR10_n, RUPT1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4015(__A04_NET_214, __A04_1__STG1, QC0_n, SQEXT_n, SQ1_n, __A04_NET_259, GND, __A04_NET_200, SUMB16_n, SUMA16_n, TSGU_n, __A04_NET_258, __A04_1__STG2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4016(__A04_NET_255, __A04_NET_258, __A04_1__ST376, DV3764, DIV_n, __A04_NET_255, GND, __A04_NET_256, __A04_1__ST376, __A04_1__ST1376_n, DIV_n, __A04_1__ST1376_n, DV1376, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U4017(__A04_NET_259, DIV_n, __A04_1__DV0, __A04_1__DV0_n, DV1, DV1_n, GND, DV376_n, __A04_1__DV376, __A04_NET_202, TL15, BR1, __A04_NET_215, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4018(__A04_1__DV0, DIV_n, ST0_n, DV1, DIV_n, ST1_n, GND, DIV_n, __A04_1__ST4_n, DV4, DIV_n, __A04_1__ST376_n, __A04_1__DV376, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4019(__A04_NET_192, SUMA16_n, SUMB16_n, __A04_NET_201, PHS4, PHS3_n, GND, UNF_n, TOV_n, __A04_NET_196, L15_n, __A04_NET_202, __A04_NET_197, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U4020(PHS4_n, WL16_n, __A04_NET_197, __A04_NET_186, __A04_NET_193, __A04_NET_185, GND, __A04_NET_184, __A04_NET_215, __A04_NET_198, __A04_NET_199, __A04_NET_186, TSGN_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4021(__A04_NET_198, TSGN_n, PHS3_n, __A04_NET_199, __A04_NET_202, PHS3_n, GND, TOV_n, PHS2_n, __A04_NET_205, __A04_1__SGUM, __A04_NET_196, __A04_NET_187, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U4022(__A04_NET_189, __A04_NET_192, PHS3_n, TSGU_n, PHS4,  , GND,  , WL16_n, WL15_n, WL14_n, WL13_n, __A04_NET_226, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U4023(__A04_NET_187, __A04_NET_215_U4023_2, __A04_NET_185, __A04_NET_215_U4023_4, __A04_NET_184, __A04_NET_193_U4023_6, GND, __A04_NET_193_U4023_8, __A04_NET_188, __A04_NET_204_U4023_10, __A04_NET_226, __A04_NET_204_U4023_12, __A04_NET_227, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U4024(__A04_NET_188, __A04_NET_205, __A04_NET_189, __A04_NET_195, TOV_n, OVF_n, GND, __A04_NET_230, PHS3_n, __A04_NET_207, TMZ_n, PHS4_n, __A04_NET_225, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U4025(__A04_NET_193, BR1_n, __A04_1__TSGN2, __A04_NET_230, __A04_NET_208, BR2, GND, BR2_n, __A04_NET_209, DV4_n, DV4, __A04_NET_281, __A04_NET_315, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4026(GEQZRO_n, PHS4_n, WL16_n, PHS4_n, __A04_NET_230, __A04_NET_203, GND, __A04_NET_211, __A04_NET_203, __A04_NET_204, __A04_NET_209, __A04_NET_194, TPZG_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U4027(__A04_NET_227, WL12_n, WL11_n, WL10_n, WL09_n,  , GND,  , WL08_n, WL07_n, WL06_n, WL05_n, __A04_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U4028(__A04_NET_223, WL04_n, WL03_n, WL02_n, WL01_n,  , GND,  , __A04_NET_208, __A04_NET_207, __A04_NET_206, __A04_NET_205, __A04_NET_209, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U4029(__A04_NET_222, __A04_NET_204_U4029_2, __A04_NET_223, __A04_NET_204_U4029_4, __A04_NET_225, __A04_NET_204_U4029_6, GND, __A04_NET_208_U4029_8, __A04_NET_210, __A04_NET_208_U4029_10, __A04_NET_211,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4030(__A04_NET_206, TMZ_n, PHS3_n, __A04_NET_210, __A04_NET_194, __A04_NET_195, GND, SQ0_n, EXST0_n, __A04_NET_315, QC3_n, SQEXT, __A04_NET_280, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4031(__A04_NET_281, SQR10, QC0_n, __A04_NET_281, SQR10_n, __A04_2__WRITE0, GND, RAND0, SQR10, __A04_NET_281, QC1_n, READ0, QC0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U4032(READ0, __A04_2__READ0_n, __A04_2__WRITE0, __A04_2__WRITE0_n, WOR0, __A04_2__WOR0_n, GND, RXOR0_n, RXOR0, __A04_2__RUPT0_n, RUPT0, __A04_2__RUPT1_n, RUPT1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4033(QC1_n, SQR10_n, SQR10, __A04_NET_281, QC2_n, ROR0, GND, WOR0, QC2_n, __A04_NET_281, SQR10_n, WAND0, __A04_NET_281, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4034(SQR10, __A04_NET_281, QC3_n, __A04_NET_281, SQR10_n, RUPT0, GND, __A04_NET_296, ST0_n, SQR12_n, SQ2_n, RXOR0, QC3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U4035(__A04_NET_296, __A04_NET_287, INOUT, INOUT_n, __A04_NET_279, __A04_NET_306, GND, BR1B2_n, __A04_2__BR1B2, BR12B_n, __A04_2__BR12B, BR1B2B_n, BR1B2B, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4036(PRINC, __A04_NET_280, __A04_NET_287, RRPA, T03_n, __A04_2__RUPT1_n, GND, T03_n, RXOR0_n, n3XP7, __A04_NET_286, T03_n, __A04_NET_283, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4037(EXST0_n, SQ0_n, INOUT, DV4, PRINC, __A04_NET_319, GND, __A04_NET_316, __A04_NET_283, __A04_NET_285, __A04_NET_275, INOUT, RUPT0, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4038(__A04_NET_286, ROR0, WOR0, __A04_NET_282, T03_n, __A04_NET_284, GND, RAND0, WAND0, __A04_NET_284, DV4_n, T05_n, n5XP28, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U4039(__A04_NET_316, RB_n_U4039_2, __A04_NET_310, RC_n_U4039_4, __A04_NET_309, n5XP11_U4039_6, GND, n5XP11_U4039_8, __A04_NET_308, RA_n_U4039_10, __A04_NET_307, WG_n_U4039_12, __A04_NET_314, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U4040(__A04_NET_282, __A04_NET_277, T05_n, INOUT_n, READ0, __A04_NET_309, GND, WCH_n, __A04_NET_276, n7XP14, __A04_NET_278, __A04_NET_310, __A04_NET_272, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4041(__A04_NET_308, __A04_2__WRITE0, RXOR0, __A04_NET_285, __A04_2__READ0_n, T05_n, GND, __A04_2__WRITE0_n, T05_n, __A04_NET_276, T05_n, __A04_2__WOR0_n, __A04_NET_278, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4042(__A04_NET_277, T05_n, RXOR0_n, __A04_NET_271, T02_n, __A04_2__WRITE0_n, GND, T02_n, INOUT_n, n2XP3, T09_n, __A04_2__RUPT0_n, n9XP1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4043(__A04_NET_276, __A04_NET_277, RUPT1, IC13, IC12, __A04_NET_273, GND, __A04_NET_314, n9XP1, __A04_NET_272, __A04_NET_275, __A04_NET_307, n2XP3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4044(__A04_NET_272, T09_n, RXOR0_n, __A04_NET_275, T09_n, __A04_NET_273, GND, __A04_NET_277, __A04_NET_271, __A04_NET_313, T01_n, __A04_2__RUPT1_n, RB2, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U4045(__A04_NET_313, WG_n_U4045_2, __A04_NET_311, __A04_NET_279_U4045_4, __A04_NET_312, __A04_NET_279_U4045_6, GND, RA_n_U4045_8, __A04_NET_327, WG_n_U4045_10, __A04_NET_329, TMZ_n_U4045_12, __A04_NET_328, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4046(RUPT0, RUPT1, INOUT, MP1, MP3A, __A04_NET_311, GND, __A04_NET_312, __A04_1__DV0, IC15, DV1376, __A04_NET_274, RSM3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4047(R15, __A04_NET_274, T01_n, n1XP10, T01_n, __A04_1__DV0_n, GND, MP0_n, T03_n, __A04_NET_299, INOUT_n, T03_n, __A04_NET_288, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4048(T02_n, __A04_1__DV0_n, BRDIF_n, TS0_n, T04_n, __A04_NET_297, GND, __A04_NET_298, T04_n, BR1, MP0_n, n2XP5, BR1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4049(n3XP2, T03_n, TS0_n, __A04_2__BR1B2, BR1, BR2_n, GND, BR1_n, BR2, __A04_2__BR12B, __A04_2__BR1B2, __A04_2__BR12B, BRDIF_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4050(BR1B2B, BR2, BR1, n4XP5, TS0_n, T04_n, GND, T04_n, INOUT_n, n4XP11, T04_n, MP3_n, __A04_NET_294, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4051(MP0_n, BR1_n, DV1_n, T04_n, BR2_n, __A04_NET_300, GND, __A04_NET_305, TS0_n, T05_n, BR1B2_n, __A04_NET_290, T04_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4052(T05_n, TS0_n, T07_n, BR1_n, MP3_n, n7XP19, GND, n8XP6, T08_n, DV1_n, BR2, __A04_NET_303, BR12B_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4053(B15X, T05_n, DV1_n, n5XP4, T05_n, RSM3_n, GND, T06_n, DV1_n, n6XP5, T06_n, MP3_n, TL15, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4054(__A04_1__TSGN2, T07_n, MP0_n, __A04_NET_301, T07_n, DV1_n, GND, T08_n, DV1_n, n8XP5, T09_n, MP3_n, __A04_NET_292, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4055(T09_n, BR1, T09_n, MP0_n, BR1_n, __A04_NET_289, GND, __A04_NET_302, MP0_n, T09_n, BRDIF_n, __A04_NET_293, MP0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4056(KRPT, T09_n, __A04_2__RUPT1_n, MP0T10, T10_n, MP0_n, GND, __A04_NET_306, T02_n, __A04_NET_295, STORE1_n, T09_n, __A04_NET_291, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U4057(BR1_n, MP0_n, n1XP10, n8XP5, __A04_NET_292, __A04_NET_327, GND, __A04_NET_337, __A04_NET_300, __A04_NET_299, __A04_NET_301, __A04_NET_304, T11_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0) U4058(DVST, __A04_1__DVST_n, __A04_NET_304, __A04_NET_336, TRSM, __A04_1__TRSM_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b1) U4059( ,  , __A04_NET_288, B15X, n7XP19, __A04_NET_323, GND, __A04_NET_322, n8XP5, __A04_NET_293, __A04_NET_289,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4060(__A04_NET_328, n2XP5, n1XP10, __A04_NET_324, __A04_NET_297, __A04_NET_302, GND, n1XP10, MP0T10, __A04_NET_325, __A04_NET_305, __A04_NET_304, __A04_NET_335, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U4061(__A04_NET_323, WY_n_U4061_2, __A04_NET_322, WY_n_U4061_4, __A04_NET_320, WL_n_U4061_6, GND, RC_n_U4061_8, __A04_NET_321, RB_n_U4061_10, __A04_NET_326, CI_n_U4061_12, __A04_NET_324, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U4062(__A04_NET_298, __A04_NET_290, __A04_NET_290, n2XP5, __A04_NET_289, __A04_NET_321, GND, __A04_NET_326, __A04_NET_298, n7XP19, __A04_NET_293, __A04_NET_320, n6XP5, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U4063(__A04_NET_325, TSGN_n_U4063_2, __A04_NET_337, TSGN_n_U4063_4, __A04_NET_335, RB1_n_U4063_6, GND, L16_n_U4063_8, __A04_NET_336, R1C_n_U4063_10, __A04_NET_334, n8PP4_U4063_12, __A04_NET_319, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U4064(__A04_NET_334, __A04_NET_304, __A04_NET_303, __A04_2__BRXP3, T03_n, IC15_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U4065(RSC_n, __A04_NET_295, __A04_NET_294, __A04_NET_301, __A04_2__BRXP3,  , GND,  , __A04_NET_295, __A04_NET_291, __A04_NET_294, __A04_2__BRXP3, __A04_NET_329, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U4066(__A04_NET_244, MST1_U4066_2, __A04_NET_257, MST2_U4066_4, __A04_NET_214, MST3_U4066_6, GND, MBR1_U4066_8, __A04_NET_215, MBR2_U4066_10, __A04_NET_208, MWCH_U4066_12, WCH_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U4067(RSC_n, MRSC_U4067_2,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U5001(IC10, IC3, TC0, TCF0, IC4, __A05_NET_217, GND, __A05_NET_215, IC2, IC3, RSM3, __A05_NET_212, IC2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5002(__A05_NET_211, STD2, IC2, __A05_NET_198, T01_n, __A05_NET_212, GND, T01_n, __A05_NET_211, __A05_NET_213, IC10_n, T01_n, __A05_NET_219, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5003(__A05_NET_218, T01_n, __A05_NET_217, __A05_NET_216, T02_n, __A05_NET_215, GND, T08_n, CCS0_n, __A05_NET_254, T02_n, MP3_n, n2XP7, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U5004(T02_n, STD2, __A05_1__10XP6, __A05_1__10XP7, __A05_NET_219, __A05_NET_214, GND, __A05_NET_209, __A05_NET_213, n3XP6, __A05_NET_188, DVST, DIV_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U5005(__A05_NET_214, MONEX_n_U5005_2, __A05_NET_209, RZ_n_U5005_4, __A05_NET_203, RB_n_U5005_6, GND, RA_n_U5005_8, __A05_NET_210, WA_n_U5005_10, __A05_NET_208, RL_n_U5005_12, __A05_NET_220, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U5006(__A05_NET_216, __A05_1__8XP15, __A05_NET_181, __A05_NET_183, __A05_1__8XP12, __A05_NET_220, GND, __A05_1__PARTC, INKL_n, SHIFT, MONpCH, NISQ_n, n2XP7, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5007(__A05_1__3XP5, T03_n, IC2_n, __A05_NET_206, T01_n, IC15_n, GND, __A05_NET_206, __A05_NET_185, __A05_NET_210, T03_n, TC0_n, n3XP6, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5008(__A05_NET_185, T04_n, IC2_n, __A05_NET_184, T02_n, IC15_n, GND, __A05_NET_184, __A05_NET_186, TPZG_n, T04_n, DAS0_n, __A05_NET_181, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U5009(__A05_NET_208, __A05_NET_181, __A05_NET_182, __A05_NET_182, T04_n, MASK0_n, GND, MP3_n, T10_n, __A05_NET_183, T05_n, IC2_n, __A05_NET_188, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5010(__A05_NET_186, T05_n, __A05_NET_187, __A05_NET_221, __A05_NET_206, __A05_NET_186, GND, T05_n, DAS0_n, n5XP12, T06_n, RSM3_n, __A05_NET_205, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U5011(__A05_1__PARTC, PRINC, __A05_NET_186, __A05_NET_206, n7XP9, __A05_NET_178, GND, __A05_NET_177, n9XP5, __A05_NET_206, __A05_NET_205, __A05_NET_187, CCS0, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U5012(__A05_NET_221, TMZ_n_U5012_2, __A05_NET_177, WG_n_U5012_4, __A05_NET_179, RG_n_U5012_6, GND, RC_n_U5012_8, __A05_NET_204, A2X_n_U5012_10, __A05_NET_193, WY_n_U5012_12, __A05_NET_189, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5013(__A05_NET_191, T06_n, DAS0_n, __A05_NET_190, T06_n, MSU0_n, GND, __A05_NET_182, __A05_NET_190, __A05_NET_204, T07_n, DAS0_n, __A05_NET_199, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b1) U5014(__A05_NET_186, __A05_NET_192, __A05_NET_192, __A05_NET_191, __A05_NET_190, __A05_NET_193, GND, __A05_NET_189, __A05_NET_192, __A05_NET_190, __A05_NET_191, __A05_NET_179, __A05_NET_191, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U5015(__A05_NET_203, __A05_NET_218, __A05_1__3XP5, __A05_NET_199, __A05_NET_205,  , GND,  , IC3, RSM3, MP3, IC16, TSUDO_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5016(n7XP9, T07_n, MSU0_n, __A05_NET_192, T07_n, IC2_n, GND, T07_n, CCS0_n, __A05_NET_248, __A05_NET_243, __A05_NET_235, __A05_NET_240, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U5017(__A05_NET_190, __A05_NET_198, __A05_1__8XP3, __A05_NET_248, n4XP5, __A05_NET_194, GND, __A05_NET_249, n4XP5, __A05_NET_248, __A05_NET_198, __A05_NET_196, __A05_1__10XP6, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U5018(__A05_NET_196, CI_n_U5018_2, __A05_NET_194, RZ_n_U5018_4, __A05_NET_249, WY12_n_U5018_6, GND, WZ_n_U5018_8, __A05_NET_244, RB_n_U5018_10, __A05_NET_240, WB_n_U5018_12, __A05_NET_246, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U5019(CCS0_n, T07_n, BR1_n, CCS0_n, T07_n, PTWOX, GND, __A05_NET_244, __A05_1__3XP5, __A05_NET_250, __A05_NET_254, n7XP4, BR2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U5020(INKL_n, FETCH0, __A05_NET_254, __A05_NET_252, n9XP5, __A05_NET_253, GND, __A05_NET_256, IC2, IC4, DXCH0, __A05_NET_243, T08_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U5021(RAD, TSUDO_n, T08_n, __A05_NET_246, RAD, __A05_NET_247, GND, T08_n, __A05_NET_245, __A05_1__8XP15, T08_n, __A05_NET_255, __A05_1__8XP3, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U5022(IC16, __A05_NET_245, __A05_NET_350, RQ_n, MP3, __A05_NET_316, GND, SCAD_n, SCAD, NDR100_n, __A05_NET_296, __A05_NET_261, __A05_NET_262, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5023(__A05_NET_255, MP0, IC1, __A05_NET_252, T08_n, __A05_NET_256, GND, T08_n, __A05_NET_257, __A05_NET_247, T08_n, GOJ1_n, RSTRT, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U5024(__A05_NET_253, RU_n_U5024_2, __A05_NET_231, RA_n_U5024_4, __A05_NET_230, ST2_n_U5024_6, GND, WY_n_U5024_8, __A05_NET_224, RC_n_U5024_10, __A05_NET_239, WA_n_U5024_12, __A05_NET_234, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U5025(DXCH0, GOJ1, CCS0_n, BR2, T10_n, __A05_1__10XP6, GND, __A05_NET_226, IC1, IC10, RUPT0, __A05_NET_257, DAS0, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5026(__A05_1__8XP12, T08_n, DAS0_n, __A05_NET_250, T08_n, TCSAJ3_n, GND, T09_n, __A05_NET_251, __A05_NET_235, IC2, __A05_1__DV1B1B, __A05_NET_251, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5027(n9XP5, T09_n, DAS0_n, __A05_NET_222, T09_n, MASK0_n, GND, __A05_NET_222, __A05_NET_223, __A05_NET_231, T10_n, CCS0_n, __A05_NET_232, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5028(__A05_NET_230, __A05_NET_250, __A05_NET_232, n10XP1, __A05_NET_226, T10_n, GND, T10_n, __A05_NET_225, __A05_NET_223, DAS0, __A05_NET_227, __A05_NET_225, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U5029(__A05_NET_232, __A05_NET_222, T10_n, DAS0_n, BR1B2_n, n10XP8, GND, __A05_NET_234, __A05_NET_235, __A05_NET_236, n5XP11, __A05_NET_224, __A05_NET_223, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5030(__A05_NET_227, MSU0_n, BR1_n, __A05_1__10XP7, T10_n, __A05_NET_228, GND, __A05_NET_227, __A05_NET_229, __A05_NET_228, BR12B_n, DAS0_n, __A05_NET_229, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5031(n11XP2, T11_n, MSU0_n, __A05_NET_237, T11_n, MASK0_n, GND, __A05_NET_222, __A05_NET_237, __A05_NET_239, T11_n, __A05_NET_238, __A05_NET_236, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5032(__A05_NET_238, MSU0, IC14, __A05_NET_293, T10_n, __A05_NET_339, GND, GOJAM, GNHNC, __A05_NET_233, __A05_NET_233, T01, GNHNC, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U5033(__A05_NET_307, __A05_NET_351, IC12, DAS0, DAS1, __A05_NET_308, GND, __A05_NET_310, RL10BB, __A05_NET_283, RSCT, __A05_NET_301, __A05_2__6XP2, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U5034( ,  ,  ,  ,  ,  , GND, __A05_NET_282_U5034_8, __A05_NET_308, __A05_NET_282_U5034_10, __A05_NET_309, WS_n_U5034_12, __A05_NET_310, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5035(__A05_2__10XP10, T10_n, IC11_n, __A05_NET_345, T10_n, __A05_NET_346, GND, T01_n, __A05_NET_282, RL10BB, T01_n, FETCH0_n, R6, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U5036(__A05_NET_309, IC9, DXCH0, PRINC, INOUT,  , GND,  , YB0_n, YT0_n, S12, S11, __A05_NET_296, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5037(__A05_NET_283, T01_n, CHINC_n, __A05_NET_349, T03_n, __A05_NET_285, GND, IC5, MP0, __A05_NET_299, T03_n, IC8_n, __A05_NET_284, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U5038(T01_n, MONpCH, TS0, DAS0, MASK0, __A05_NET_302, GND, __A05_NET_300, __A05_NET_349, __A05_NET_284, __A05_NET_350, RSCT, INKL_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U5039(__A05_NET_300, WB_n_U5039_2, __A05_NET_301, WB_n_U5039_4, __A05_NET_302, __A05_NET_285_U5039_6, GND, __A05_NET_285_U5039_8, __A05_NET_299, RL_n_U5039_10, __A05_NET_298, RA_n_U5039_12, __A05_NET_303, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5040(n2XP8, T02_n, FETCH0_n, __A05_NET_350, T03_n, QXCH0_n, GND, T04_n, DV1_n, __A05_NET_305, T04_n, __A05_NET_306, __A05_NET_307, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U5041(__A05_NET_284, __A05_NET_305, DV1, INOUT, IC2, __A05_NET_306, GND, __A05_NET_327, __A05_NET_351, __A05_NET_348, __A05_2__5XP9, __A05_NET_298, __A05_2__11XP6, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5042(__A05_NET_303, __A05_NET_349, __A05_2__6XP2, TRSM, T05_n, NDX0_n, GND, IC12_n, T05_n, __A05_NET_351, DAS1_n, T05_n, __A05_NET_348, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U5043(__A05_2__5XP13, n5XP15, DAS1, PRINC, __A05_1__PARTC, __A05_NET_325, GND, __A05_NET_326, __A05_NET_328, n2XP8, __A05_2__10XP10, __A05_NET_324, __A05_NET_318, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U5044(__A05_NET_327, RG_n_U5044_2, __A05_NET_324, RG_n_U5044_4, __A05_NET_326, WY_n_U5044_6, GND, A2X_n_U5044_8, __A05_NET_333, CI_n_U5044_10, __A05_NET_330, WY12_n_U5044_12, __A05_NET_313, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U5045(__A05_NET_328, __A05_NET_325, T05_n, __A05_NET_333, __A05_NET_348, __A05_2__10XP10, GND, SHIFT_n, T05_n, __A05_2__5XP9, SHANC_n, T05_n, __A05_NET_331, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U5046(__A05_NET_331, __A05_NET_314, YT0_n, YB0_n, XT0_n, __A05_NET_319, GND, __A05_NET_279, RAND0, WAND0, __A05_NET_262, __A05_NET_330, __A05_NET_315, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5047(__A05_2__5XP13, IC8_n, T05_n, n5XP15, QXCH0_n, T05_n, GND, CHINC_n, T05_n, n5XP21, IC5_n, T05_n, __A05_NET_318, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U5048(__A05_NET_314, IC16_n, T05_n, __A05_NET_315, __A05_NET_316, T05_n, GND, __A05_NET_314, __A05_NET_315, __A05_NET_313, S11, S12, __A05_NET_320, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U5049(__A05_NET_317, RB_n_U5049_2, __A05_NET_323, RZ_n_U5049_4, __A05_NET_320, SCAD_U5049_6, GND, SCAD_U5049_8, __A05_NET_319, RC_n_U5049_10, __A05_NET_276, __A05_NET_260_U5049_12, __A05_NET_258, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5050(__A05_NET_317, __A05_2__5XP19, __A05_NET_314, __A05_NET_323, __A05_2__6XP7, __A05_NET_315, GND, XT2_n, NDR100_n, OCTAD2, NDR100_n, XT3_n, OCTAD3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5051(OCTAD4, NDR100_n, XT4_n, OCTAD5, NDR100_n, XT5_n, GND, NDR100_n, XT6_n, OCTAD6, BR1_n, DV1_n, __A05_NET_262, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5052(__A05_NET_280, __A05_NET_279, T05_n, __A05_2__5XP19, T05_n, __A05_NET_272, GND, DV1_n, BR1, __A05_1__DV1B1B, TS0_n, BRDIF_n, __A05_NET_264, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U5053(__A05_NET_276, __A05_NET_280, __A05_NET_281, __A05_NET_277, __A05_NET_273,  , GND,  , __A05_2__5XP13, __A05_NET_287, __A05_NET_338, __A05_NET_345, __A05_NET_335, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U5054(ROR0, __A05_1__DV1B1B, IC2, IC5, READ0, __A05_NET_258, GND, __A05_NET_265, IC2, IC3, TS0, __A05_NET_272, WOR0, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U5055(__A05_NET_259, __A05_NET_264, DV4, __A05_NET_270, __A05_NET_260, T05_n, GND, __A05_NET_261, T05_n, __A05_NET_263, __A05_NET_270, __A05_NET_281, __A05_NET_271, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U5056(__A05_NET_259, __A05_NET_260_U5056_2, __A05_NET_269, Z16_n_U5056_4, __A05_NET_271, WA_n_U5056_6, GND, __A05_NET_267_U5056_8, __A05_NET_265, __A05_NET_267_U5056_10, __A05_NET_266, WZ_n_U5056_12, __A05_NET_268, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0) U5057(__A05_NET_263, __A05_NET_269, __A05_NET_352, __A05_NET_268, __A05_NET_281, __A05_NET_341, GND, __A05_NET_334, __A05_NET_277, NISQ, NISQ_n,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U5058(__A05_NET_266, IC16, MP3, __A05_NET_352, T06_n, __A05_NET_267, GND, T06_n, DAS1_n, n6XP8, n6XP8, __A05_2__6XP7, __A05_NET_289, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U5059(__A05_NET_289, TOV_n_U5059_2, __A05_NET_286, RU_n_U5059_4, __A05_NET_288, RU_n_U5059_6, GND, WB_n_U5059_8, __A05_NET_291, RG_n_U5059_10, __A05_NET_292, TSGN_n_U5059_12, __A05_NET_342, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5060(__A05_2__6XP7, DV4_n, T06_n, __A05_NET_340, T07_n, __A05_NET_297, GND, T07_n, STFET1_n, __A05_NET_294, T08_n, DV4_n, RSTSTG, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U5061(__A05_NET_352, n6XP8, __A05_NET_293, __A05_NET_338, __A05_NET_287, __A05_NET_288, GND, __A05_2__6XP2, T06_n, RXOR0, INOUT_n, __A05_NET_286, n5XP11, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U5062(IC13, IC14, __A05_NET_340, __A05_NET_338, __A05_NET_293, __A05_NET_291, GND, __A05_NET_292, __A05_NET_340, __A05_NET_294, __A05_NET_273, __A05_NET_297, DV1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U5063(T08_n, MONWBK, IC2, IC14, DV1, __A05_NET_339, GND, __A05_NET_346, DV4B1B, IC4, __A05_NET_344, U2BBK, STFET1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U5064(__A05_NET_342, RSTSTG, __A05_2__5XP9, __A05_NET_281, T09_n, __A05_NET_261, GND, T09_n, DV4_n, __A05_NET_338, T09_n, DAS1_n, __A05_NET_277, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U5065(__A05_NET_341, Z15_n_U5065_2, __A05_NET_335, WL_n_U5065_4, __A05_NET_334, TMZ_n_U5065_6, GND, WYD_n_U5065_8, __A05_NET_343, TSGN_n_U5065_10, __A05_NET_178,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U5066(DAS1_n, ADS0, T12_n, T12USE_n, DV1_n, __A05_NET_287, GND,  ,  ,  ,  , __A05_NET_344, BR2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U5067(DV4B1B, DV4_n, BR1, __A05_2__11XP6, T11_n, DV1_n, GND, __A05_2__5XP9, __A05_2__11XP6, __A05_NET_343, T11_n, RXOR0_n, __A05_NET_273, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U5068(NISQ_n, MNISQ_U5068_2,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U6001(T04, T07, __A06_NET_273, __A06_NET_309, __A06_NET_271, __A06_NET_275, GND, __A06_NET_308, T01, T03, T05, __A06_NET_274, T10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6002(__A06_NET_273, __A06_NET_274, DV376_n, __A06_NET_309, T01_n, DV1376_n, GND, T04_n, DV4_n, __A06_NET_271, MP1_n, __A06_NET_272, __A06_NET_276, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U6003(T07, T09, __A06_NET_288, __A06_1__L02A_n, L01_n, __A06_NET_292, GND, __A06_NET_352, T05, T08, T11, __A06_NET_310, T11, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U6004(__A06_NET_308, __A06_NET_272_U6004_2, __A06_NET_310, __A06_NET_272_U6004_4, __A06_NET_304, A2X_n_U6004_6, GND, RB_n_U6004_8, __A06_NET_307, WYD_n_U6004_10, __A06_NET_306, WY_n_U6004_12, __A06_NET_322, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0) U6005(__A06_NET_321, __A06_NET_276, n2XP7, L2GD_n, __A06_1__ZIP, __A06_1__DVXP1, GND, __A06_1__DVXP1, __A06_NET_300, __A06_NET_306, __A06_NET_302, __A06_NET_303, __A06_NET_301, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U6006(L01_n, __A06_NET_299, __A06_1__L02A_n, __A06_NET_289, __A06_NET_288, __A06_NET_305, GND, __A06_1__DVXP1, __A06_NET_275, __A06_1__ZIP, __A06_NET_321, __A06_NET_293, __A06_NET_291, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U6007(n7XP19, __A06_1__ZIP, __A06_1__DVXP1, __A06_NET_290, RBSQ, __A06_NET_307, GND, __A06_NET_298, __A06_NET_299, __A06_NET_289, __A06_NET_305, __A06_NET_304, __A06_1__DVXP1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U6008(__A06_NET_305, __A06_NET_299, __A06_NET_321, __A06_NET_303, __A06_NET_302, __A06_NET_323, GND, __A06_NET_291, __A06_NET_302, __A06_NET_303, __A06_1__L02A_n, __A06_NET_303, __A06_1__L02A_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6009(__A06_NET_300, __A06_NET_321, __A06_NET_301, __A06_NET_294, __A06_NET_321, __A06_NET_293, GND, __A06_NET_352, DV376_n, __A06_NET_297, DV1376_n, T02_n, __A06_NET_296, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U6010(__A06_NET_294, MCRO_n, __A06_NET_295, __A06_NET_346, __A06_NET_313, __A06_NET_287, GND, __A06_1__ZAP, ZAP_n, __A06_NET_348, __A06_NET_352, MONEX, MONEX_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U6011(__A06_NET_321, __A06_NET_293, __A06_NET_291, __A06_NET_298, __A06_NET_321, __A06_NET_290, GND, __A06_NET_302, __A06_NET_289, __A06_NET_288, L01_n, __A06_1__ZIPCI, __A06_NET_292, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0) U6012(__A06_NET_295, __A06_NET_297, __A06_NET_296, __A06_NET_313, __A06_NET_314, DIVSTG, GND, T08, T10, __A06_NET_311, MP1_n, __A06_NET_320, __A06_NET_319, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U6013(T06, T09, DV376_n, __A06_NET_315, T12USE_n, __A06_NET_314, GND, __A06_NET_312, T02, T04, T06, __A06_NET_315, T12, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U6014(__A06_NET_312, __A06_NET_320_U6014_2, __A06_NET_311, __A06_NET_320_U6014_4, __A06_NET_316, WL_n_U6014_6, GND, RG_n_U6014_8, __A06_NET_280, WB_n_U6014_10, __A06_NET_277, RU_n_U6014_12, __A06_NET_284, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U6015(__A06_NET_318, T01, T03, __A06_NET_317, __A06_NET_318, MP3_n, GND, __A06_NET_319, __A06_NET_317, ZAP_n, n5XP28, __A06_NET_346, TSGU_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b1) U6016(__A06_NET_316, __A06_NET_346, n5XP12, __A06_NET_283, RRPA, n5XP4, GND, n5XP15, n3XP6, WQ_n, n9XP5, n6XP8, __A06_NET_351, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U6017(__A06_NET_280, n5XP4, RADRG, __A06_NET_346, n5XP28,  , GND,  , n5XP28, n1XP10, __A06_NET_287, n2XP3, __A06_NET_277, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U6018(__A06_NET_284, __A06_NET_287, __A06_1__ZAP, n5XP12, n6XP5,  , GND,  , PRINC, PINC, MINC, DINC, __A06_NET_258, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U6019(__A06_NET_283, WZ_n_U6019_2, __A06_NET_345, TOV_n_U6019_4, __A06_NET_351, WSC_n_U6019_6, GND, WG_n_U6019_8, __A06_NET_350, __A06_NET_203_U6019_10, __A06_NET_270, __A06_NET_203_U6019_12, __A06_NET_236, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U6020(n6XP5, n3XP2, BR1_n, PHS4_n, TSGU_n, RB1F, GND, CLXC, TSGU_n, BR1, PHS4_n, __A06_NET_345, n9XP5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b1) U6021(__A06_NET_350, n6XP8, n6XP8, PIFL_n, __A06_1__DVXP1, __A06_NET_347, GND, PTWOX, MONEX, __A06_NET_332, MONEX, B15X, __A06_NET_331, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U6022(PIFL_n, __A06_NET_348, STBE, n1XP10, STBF, __A06_NET_326, GND, __A06_NET_270, __A06_NET_205, __A06_NET_206, INCR0, __A06_NET_347, T02, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0) U6023(__A06_NET_332, TWOX, __A06_NET_331, BXVX, __A06_NET_333, __A06_NET_336, GND, __A06_NET_335, __A06_NET_336, __A06_NET_334, __A06_NET_335, __A06_NET_327, __A06_NET_334, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U6024(CGMC, __A06_NET_326, __A06_NET_324, __A06_NET_337, CGMC, __A06_NET_333, GND, __A06_NET_337, __A06_NET_326, __A06_NET_333, BR1, AUG0_n, __A06_NET_205, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0) U6025(__A06_NET_327, __A06_NET_328, __A06_NET_328, __A06_NET_330, __A06_NET_330, __A06_NET_329, GND, __A06_NET_324, __A06_NET_329, __A06_NET_240, __A06_NET_242, __A06_NET_253, __A06_2__7XP10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6026(__A06_NET_206, DIM0_n, BR12B_n, __A06_NET_236, PINC, __A06_NET_204, GND, BR12B_n, DINC_n, __A06_NET_204, T06_n, __A06_NET_203, __A06_2__6XP10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6027(__A06_NET_231, MINC, MCDU, __A06_NET_234, AUG0_n, BR1_n, GND, DIM0_n, BR1B2B_n, __A06_NET_233, BR1B2B_n, DINC_n, __A06_NET_232, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U6028(__A06_NET_234, __A06_NET_233, BR1B2B_n, CDUSTB_n, DINC_n, __A06_2__POUT, GND, __A06_2__MOUT, BR12B_n, CDUSTB_n, DINC_n, __A06_NET_230, __A06_NET_232, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U6029(__A06_NET_231, __A06_NET_241_U6029_2, __A06_NET_230, __A06_NET_241_U6029_4, __A06_NET_240, MONEX_n_U6029_6, GND, WA_n_U6029_8, __A06_NET_222, RB1_n_U6029_10, __A06_NET_253, R1C_n_U6029_12, __A06_NET_250, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6030(__A06_NET_242, T06_n, __A06_NET_241, __A06_NET_239, PCDU, MCDU, GND, T06_n, __A06_NET_239, __A06_2__6XP12, __A06_NET_224, T07_n, __A06_NET_223, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b1) U6031(BR2_n, DINC_n, DAS0, DAS1, MSU0, __A06_NET_224, GND, __A06_NET_222, __A06_NET_223, __A06_2__7XP7, __A06_NET_221, __A06_2__ZOUT, CDUSTB_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6032(__A06_NET_229, DV4_n, BR1B2B, __A06_2__7XP7, T07_n, __A06_NET_228, GND, WAND0, INOTLD, __A06_NET_226, T07_n, __A06_NET_226, n7XP14, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U6033(__A06_NET_229, WAND0, DAS1_n, T07_n, BR1B2_n, __A06_2__7XP10, GND, __A06_2__7XP11, DAS1_n, T07_n, BR12B_n, __A06_NET_228, RAND0, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U6034(__A06_2__7XP11, __A06_NET_250, __A06_NET_191, PONEX, ST2_n, ST2, GND, ST1, __A06_NET_207, __A06_NET_267, PSEUDO, __A06_NET_266, __A06_2__RDBANK, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6035(__A06_2__7XP15, __A06_NET_251, T07_n, __A06_NET_257, __A06_NET_258, T07_n, GND, PRINC, INKL, __A06_NET_246, IC9, DXCH0, __A06_NET_249, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U6036(PCDU, MCDU, n7XP9, n11XP2, __A06_2__7XP15, RUS_n, GND, __A06_NET_255, __A06_NET_257, __A06_NET_256, __A06_NET_221, __A06_NET_251, SHIFT, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U6037(__A06_NET_255, RU_n_U6037_2, __A06_NET_243, WSC_n_U6037_4, __A06_NET_245, WG_n_U6037_6, GND, RB_n_U6037_8, __A06_NET_248, n8PP4_U6037_10, __A06_NET_247, n8PP4_U6037_12, __A06_NET_196, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U6038(__A06_NET_246, T07_n, T04_n, MON_n, FETCH1, __A06_NET_244, GND, __A06_NET_243, __A06_NET_269, __A06_NET_244, __A06_NET_268, __A06_NET_269, MONpCH, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6039(__A06_NET_245, __A06_NET_269, __A06_NET_268, __A06_NET_268, T07_n, __A06_NET_249, GND, __A06_2__10XP9, __A06_NET_268, __A06_NET_248, T08_n, n8PP4, __A06_2__8XP4, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U6040(RUPT1, DAS1, IC17, MASK0, IC11, __A06_NET_196, GND, __A06_NET_195, IC6, IC7, IC9, __A06_NET_247, MSU0, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U6041(__A06_NET_195, n8PP4_U6041_2, __A06_NET_193, __A06_NET_199_U6041_4, __A06_NET_192, __A06_NET_199_U6041_6, GND, WS_n_U6041_8, __A06_NET_197, __A06_NET_186_U6041_10, __A06_NET_185, __A06_NET_186_U6041_12, __A06_NET_184, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U6042(T08_n, RUPT0, __A06_NET_199, R6, R15, __A06_NET_197, GND, __A06_NET_184, ADS0, IC11, __A06_NET_183, __A06_NET_193, DAS0, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6043(__A06_NET_192, MP1, DV1376, __A06_NET_198, MP3_n, BR1_n, GND, __A06_NET_198, CCS0, __A06_NET_185, T11_n, __A06_NET_186, __A06_NET_221, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6044(__A06_NET_183, DAS1_n, BR2_n, __A06_NET_190, __A06_1__ZIPCI, __A06_2__6XP12, GND, CCS0_n, BR1B2B_n, __A06_NET_217, T10_n, NDXX1_n, EXT, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U6045(T03_n, DAS1_n, __A06_NET_209, __A06_NET_256, n2XP5, __A06_NET_208, GND, __A06_NET_216, IC7, DCS0, SU0, __A06_NET_256, ADS0, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U6046(__A06_NET_191, n8XP6, n7XP4, n10XP8, __A06_2__6XP10,  , GND,  , IC6, DCA0, AD0, __A06_NET_217, __A06_NET_211, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U6047(__A06_NET_190, CI_n_U6047_2, __A06_NET_208, WA_n_U6047_4, __A06_NET_213, RC_n_U6047_6, GND, __A06_NET_220_U6047_8, __A06_NET_216, __A06_NET_220_U6047_10, __A06_NET_215, ST2_n_U6047_12, __A06_NET_200, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6048(__A06_2__10XP9, T10_n, __A06_NET_211, __A06_NET_210, IC6, IC7, GND, T10_n, __A06_NET_210, __A06_NET_209, T10_n, __A06_NET_220, __A06_NET_219, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U6049(__A06_NET_213, __A06_NET_219, __A06_2__7XP7, __A06_NET_215, __A06_NET_214, DV4B1B, GND, CCS0_n, BR12B_n, __A06_NET_214, T10_n, MP1_n, __A06_2__10XP15, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U6050(__A06_2__8XP4, __A06_2__10XP15, __A06_2__8XP4, RADRZ, n9XP1, __A06_NET_264, GND, NEAC, __A06_NET_262, TL15, GOJAM, __A06_NET_200, RADRZ, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U6051(__A06_NET_207, n2XP8, n10XP1, MP0T10, __A06_2__10XP15,  , GND,  , __A06_1__DVXP1, GOJAM, NISQ, __A06_1__WHOMP_n, WHOMP, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U6052(__A06_NET_264, RZ_n_U6052_2, __A06_NET_267, RPTSET_U6052_4, __A06_NET_266, RU_n_U6052_6, GND, RC_n_U6052_8, __A06_NET_325,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U6053(__A06_NET_262, MP0T10, NEAC, __A06_NET_265, RADRZ, PSEUDO, GND, T06_n, STFET1_n, __A06_2__RDBANK, __A06_1__ZIPCI, n3XP7, __A06_NET_325, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U6054(__A06_NET_265, GOJAM, n3XP7, n5XP21, n4XP11, RCH_n, GND,  ,  ,  ,  , PSEUDO, RADRG, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U6055(R1C_n, R1C, RB1_n, RB1, L02_n, __A06_NET_341, GND, __A06_1__L02A_n, __A06_NET_341, __A06_NET_339, L15_n, __A06_NET_288, __A06_NET_339, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U6056(__A06_NET_323, __A06_NET_322, __A06_1__WHOMP_n, WHOMPA, __A06_NET_269, WOVR_n, GND, POUT_n, __A06_2__POUT, MOUT_n, __A06_2__MOUT, ZOUT_n, __A06_2__ZOUT, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U6057(__A06_1__WHOMP_n, WHOMP, CLXC,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U6058(RCH_n, MRCH_U6058_2,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U7001(__A07_1__WALSG, ZAP_n, WT_n, __A07_NET_159, __A07_NET_150, __A07_NET_160, GND, __A07_NET_159, WT_n, __A07_NET_162, WY_n, WT_n, __A07_NET_164, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0) U7002(__A07_1__WALSG, WALSG_n, WY12_n, __A07_NET_150, WY_n, __A07_NET_160, GND, WYLOG_n, __A07_NET_162, WYHIG_n, __A07_NET_164,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U7003(__A07_NET_161, __A07_NET_162, __A07_NET_163, __A07_NET_163, WYD_n, WT_n, GND, __A07_NET_161, CT_n, CUG, L15_n, PIFL_n, __A07_NET_156, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1) U7004(__A07_NET_163, WYDG_n, __A07_NET_158, WYDLOG_n, __A07_NET_157, WBG_n, GND,  ,  ,  ,  , WG1G_n, __A07_1__WGNORM, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U7005(__A07_NET_154, WYD_n, WT_n, __A07_NET_157, WB_n, WT_n, GND, WBG_n, CT_n, CBG, __A07_1__WGNORM, __A07_NET_171, WG2G_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U7006(SHIFT, NEAC, __A07_1__WGA_n, WT_n, GINH, __A07_1__WGNORM, GND, __A07_NET_171, __A07_1__WGA_n, WT_n, SR_n, __A07_NET_155, __A07_NET_156, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U7007(__A07_NET_154, __A07_NET_158_U7007_2, __A07_NET_155, __A07_NET_158_U7007_4,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U7008(__A07_1__WGA_n, WT_n, __A07_1__WGA_n, WT_n, CYL_n, __A07_NET_167, GND, __A07_NET_165, __A07_1__WGA_n, WT_n, EDOP_n, __A07_NET_170, CYR_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0) U7009(__A07_NET_170, WG5G_n, __A07_NET_167, WG3G_n, __A07_NET_165, WEDOPG_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U7010(WG4G_n, __A07_NET_171, __A07_NET_170, __A07_NET_166, WT_n, WZ_n, GND, __A07_1__WSCG_n, XB5_n, __A07_NET_168, __A07_NET_166, __A07_NET_168, WZG_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U7011(CZG, WZG_n, CT_n, __A07_NET_140, WL_n, WT_n, GND, __A07_1__WSCG_n, XB1_n, __A07_NET_143, __A07_NET_135, CT_n, CLG1G, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U7012(XB1_n, XT0_n, __A07_NET_140, __A07_NET_139, __A07_NET_143, WLG_n, GND, __A07_NET_137, __A07_NET_133, __A07_NET_138, __A07_1__WALSG, __A07_NET_139, WCHG_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U7013(__A07_NET_134, __A07_NET_140, __A07_NET_139, __A07_NET_143, __A07_1__WALSG,  , GND,  , __A07_NET_143, __A07_NET_139, __A07_NET_140, __A07_2__G2LSG, __A07_NET_135, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U7014(CLG2G, __A07_NET_134, CT_n, __A07_NET_133, WT_n, WA_n, GND, __A07_1__WSCG_n, XB0_n, __A07_NET_138, __A07_NET_133, __A07_NET_138, WAG_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U7015(CAG, __A07_NET_137, CT_n, __A07_NET_136, WT_n, WS_n, GND, WSG_n, CT_n, CSG, WT_n, WQ_n, __A07_NET_152, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1) U7016(__A07_NET_136, WSG_n,  ,  ,  ,  , GND,  ,  , RCG_n, __A07_NET_206, G2LSG_n, __A07_2__G2LSG, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U7017(__A07_NET_152, __A07_NET_151, XB2_n, XT0_n, WCHG_n, __A07_NET_153, GND,  ,  ,  ,  , WQG_n, __A07_NET_153, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U7018(__A07_NET_151, __A07_1__WSCG_n, XB2_n, CQG, WQG_n, CT_n, GND, RT_n, RC_n, __A07_NET_206, RT_n, RQ_n, __A07_NET_207, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U7019(__A07_NET_207, __A07_NET_201, XB2_n, XT0_n, RCHG_n, __A07_NET_202, GND, RFBG_n, __A07_NET_203, __A07_NET_204, __A07_2__RBBK, RQG_n, __A07_NET_202, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U7020(__A07_NET_201, __A07_2__RSCG_n, XB2_n, __A07_NET_203, __A07_2__RSCG_n, XB4_n, GND, __A07_2__RSCG_n, XB6_n, __A07_NET_204, __A07_NET_204, __A07_2__RBBK, RBBEG_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U7021(__A07_2__G2LSG, TT_n, ZAP_n, __A07_NET_208, TT_n, L2GD_n, GND, TT_n, A2X_n, __A07_NET_209, T10_n, STFET1_n, __A07_2__RBBK, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1) U7022(__A07_NET_208, L2GDG_n, __A07_NET_209, A2XG_n, __A07_NET_199, CGG, GND,  ,  ,  ,  , WBBEG_n, __A07_NET_200, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U7023(__A07_NET_197, L2GD_n, CT_n, __A07_NET_198, CT_n, WG_n, GND, __A07_1__WSCG_n, XB3_n, __A07_NET_194, __A07_NET_195, CT_n, CEBG, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U7024(__A07_NET_197, __A07_NET_198, __A07_NET_194, U2BBK, __A07_NET_200, __A07_NET_195, GND, __A07_NET_196, __A07_NET_200, U2BBK, __A07_NET_210, __A07_NET_199, CGMC, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U7025(CFBG, __A07_NET_196, CT_n, __A07_NET_210, __A07_1__WSCG_n, XB4_n, GND, __A07_NET_210, __A07_NET_200, WFBG_n, __A07_1__WSCG_n, XB6_n, __A07_NET_200, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U7026( ,  , __A07_NET_180, RGG_n,  ,  , GND,  ,  ,  ,  , REBG_n, __A07_NET_172, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U7027(__A07_NET_180, RT_n, RG_n, __A07_NET_178, RT_n, RA_n, GND, __A07_NET_178, __A07_NET_179, RAG_n, XB0_n, __A07_2__RSCG_n, __A07_NET_179, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U7028(__A07_NET_182, RT_n, RL_n, __A07_NET_183, __A07_2__RSCG_n, XB1_n, GND, RT_n, RZ_n, __A07_NET_174, __A07_NET_174, __A07_NET_173, RZG_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U7029(__A07_NET_182, __A07_NET_183, XB1_n, XT0_n, RCHG_n, __A07_NET_181, GND, US2SG, __A07_2__RUSG_n, SUMA15_n, SUMB15_n, RLG_n, __A07_NET_181, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U7030(__A07_NET_173, XB5_n, __A07_2__RSCG_n, __A07_NET_172, __A07_2__RSCG_n, XB3_n, GND, RT_n, RU_n, __A07_NET_177, RT_n, RUS_n, __A07_NET_176, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U7031(__A07_NET_177, RUG_n, __A07_NET_176, __A07_2__RUSG_n,  ,  , GND, RBHG_n, __A07_NET_191, __A07_NET_187, RL10BB,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U7032(RULOG_n, __A07_NET_177, __A07_NET_176, __A07_NET_191, RT_n, RB_n, GND, RT_n, __A07_NET_187, __A07_NET_188, __A07_NET_191, __A07_NET_188, RBLG_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0) U7033(__A07_NET_194, WEBG_n,  ,  ,  ,  , GND, __A07_NET_190, CI_n, __A07_1__WSCG_n, __A07_NET_148, __A07_2__RSCG_n, __A07_NET_186, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U7034( ,  , NEAC, EAC_n, MP3A, __A07_2__CINORM, GND, __A07_NET_186, RT_n, RSC_n, SCAD_n,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U7035(__A07_NET_189, __A07_NET_190, __A07_2__CIFF, __A07_2__CIFF, __A07_NET_189, CUG, GND, __A07_2__CIFF, __A07_2__CINORM, CI01_n, WSC_n, SCAD_n, __A07_NET_148, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U7036(__A07_NET_184, RT_n, RCH_n, __A07_NET_146, WT_n, WCH_n, GND, WCH_n, CT_n, __A07_NET_147,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1) U7037(__A07_NET_184, RCHG_n, __A07_NET_146, WCHG_n, __A07_NET_147, CCHG_n, GND, __A07_NET_149, WG_n, __A07_1__WGA_n, __A07_NET_149, U2BBKG_n, U2BBK, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U7038(__A07_NET_161, MWYG_U7038_2, WBG_n, MWBG_U7038_4, __A07_1__WGA_n, MWG_U7038_6, GND, MWZG_U7038_8, WZG_n, MWLG_U7038_10, WLG_n, MWAG_U7038_12, WAG_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U7039(WSG_n, MWSG_U7039_2, WQG_n, MWQG_U7039_4, WEBG_n, MWEBG_U7039_6, GND, MWFBG_U7039_8, WFBG_n, MWBBEG_U7039_10, WBBEG_n, MRGG_U7039_12, RGG_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U7040(RAG_n, MRAG_U7040_2, RLG_n, MRLG_U7040_4, RULOG_n, MRULOG_U7040_6, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8001(__A08_NET_203, A2XG_n, __A08_1___A1_n, __A08_NET_205, WYLOG_n, WL01_n, GND, WL16_n, WYDLOG_n, __A08_NET_198, __A08_1__Y1_n, CUG, __A08_1__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8002(PONEX, __A08_NET_203, __A08_1__X1_n, CLXC, CUG, __A08_1__X1, GND, __A08_1__Y1_n, __A08_NET_205, __A08_NET_198, __A08_1__Y1, __A08_1__X1_n, __A08_1__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8003(__A08_NET_209, __A08_1__X1_n, __A08_1__Y1_n, XUY01_n, __A08_1__X1, __A08_1__Y1, GND, __A08_NET_209, XUY01_n, __A08_NET_207, __A08_NET_209, SUMA01_n, __A08_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8004(__A08_NET_277, __A08_NET_276, SUMA01_n, SUMB01_n, RULOG_n, __A08_NET_186, GND, __A08_NET_190, __XUY03_n, XUY01_n, CI01_n, __A08_NET_278, __A08_NET_255, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U8005(CI01_n, __A08_NET_206, G01_n, GEM01, RL01_n, WL01, GND, WL01_n, WL01,  ,  , __A08_NET_154, __A08_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8006(SUMB01_n, __A08_NET_207, __A08_NET_206, __A08_NET_189, WAG_n, WL01_n, GND, WL03_n, WALSG_n, __A08_NET_191, __A08_1___A1_n, CAG, __A08_NET_187, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8007(__A08_NET_190, __CO04_U8007_2, __A08_NET_185, RL01_n_U8007_4, __A08_NET_194, L01_n_U8007_6, GND, __A08_1___Z1_n_U8007_8, __A08_NET_221, RL01_n_U8007_10, __A08_NET_220, RL01_n_U8007_12, __A08_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8008(__A08_NET_184, RAG_n, __A08_1___A1_n, __A08_NET_188, WLG_n, WL01_n, GND, __G04_n, G2LSG_n, __A08_NET_196, L01_n, CLG1G, __A08_NET_197, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8009(__A08_NET_274, WG1G_n, WL04_n, __A08_NET_193, WQG_n, WL01_n, GND, __A08_NET_193, __A08_NET_192, __A08_1___Q1_n, __A08_1___Q1_n, CQG, __A08_NET_192, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8010(__A08_NET_195, RQG_n, __A08_1___Q1_n, __A08_NET_223, WZG_n, WL01_n, GND, __A08_NET_223, __A08_NET_224, __A08_NET_221, __A08_1___Z1_n, CZG, __A08_NET_224, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8011(__A08_1___RL_OUT_1, __A08_NET_195, MDT01, RB1, R15, __A08_NET_222, GND, __A08_NET_227, __A08_NET_226, __A08_NET_225, __A08_NET_210, __A08_NET_220, __A08_NET_219, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8012(__A08_NET_219, RZG_n, __A08_1___Z1_n, __A08_NET_228, WBG_n, WL01_n, GND, __A08_NET_228, __A08_NET_229, __A08_1___B1_n, __A08_1___B1_n, CBG, __A08_NET_229, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8013(__A08_NET_171, __CO04_U8013_2, __A08_NET_227, RL01_n_U8013_4, __A08_NET_215, G01_n_U8013_6, GND, G01_n_U8013_8, __A08_NET_218, RL02_n_U8013_10, __A08_NET_142, L02_n_U8013_12, __A08_NET_143, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8014(__A08_NET_226, RBLG_n, __A08_1___B1_n, __A08_NET_225, __A08_NET_229, RCG_n, GND, WL16_n, WG3G_n, __A08_NET_214, WL02_n, WG4G_n, __A08_NET_213, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8015(__A08_NET_189, __A08_NET_191, __A08_NET_186, __A08_NET_184, CH01, __A08_NET_185, GND, __A08_NET_194, __A08_NET_188, __A08_NET_196, __A08_NET_197, __A08_1___A1_n, __A08_NET_187, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8016(__A08_NET_217, L2GDG_n, MCRO_n, __A08_NET_216, WG1G_n, WL01_n, GND, G01_n, CGG, G01, RGG_n, G01_n, __A08_NET_210, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U8017(__A08_NET_217, __A08_NET_216, WHOMPA, __XUY04_n, XUY02_n, __A08_NET_171, GND, __A08_1___RL_OUT_1, RLG_n, L01_n, GND, __A08_NET_218, G01, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U8018(__A08_NET_215, G01ED, SA01, __A08_NET_214, __A08_NET_213,  , GND,  , G02ED, SA02, __A08_NET_165, __A08_NET_164, __A08_NET_163, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8019(__A08_NET_156, A2XG_n, __A08_1___A2_n, __A08_NET_160, WYLOG_n, WL02_n, GND, WL01_n, WYDG_n, __A08_NET_159, __A08_1__Y2_n, CUG, __A08_1__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8020(TWOX, __A08_NET_156, __A08_1__X2_n, CLXC, CUG, __A08_1__X2, GND, __A08_1__Y2_n, __A08_NET_160, __A08_NET_159, __A08_1__Y2, __A08_1__X2_n, __A08_1__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8021(__A08_NET_155, __A08_1__X2_n, __A08_1__Y2_n, XUY02_n, __A08_1__X2, __A08_1__Y2, GND, __G04_n, CGG, G04, __A08_NET_155, XUY02_n, __A08_NET_150, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U8022(__A08_NET_272, __A08_NET_274, __A08_NET_155, SUMA02_n, GND, __CI03_n, GND, __A08_NET_204, SUMA02_n, SUMB02_n, RULOG_n, __A08_NET_273, G04, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8023(SUMB02_n, __A08_NET_150, __A08_NET_154, __A08_NET_157, WAG_n, WL02_n, GND, WL04_n, WALSG_n, __A08_NET_158, __A08_1___A2_n, CAG, __A08_NET_141, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8024(__A08_NET_157, __A08_NET_158, __A08_NET_204, __A08_NET_140, CH02, __A08_NET_142, GND, __A08_NET_143, __A08_NET_175, __A08_NET_172, __A08_NET_176, __A08_1___A2_n, __A08_NET_141, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8025(__A08_NET_140, RAG_n, __A08_1___A2_n, __A08_NET_175, WLG_n, WL02_n, GND, G05_n, G2LSG_n, __A08_NET_172, L02_n, CLG1G, __A08_NET_176, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8026(RLG_n, L02_n, __A08_1___RL_OUT_2, __A08_NET_144, __A08_NET_147, __A08_NET_137, GND, __A08_NET_139, MDT02, R1C, RB2, __A08_1___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8027(__A08_NET_174, WQG_n, WL02_n, __A08_1___Q2_n, __A08_NET_174, __A08_NET_146, GND, __A08_1___Q2_n, CQG, __A08_NET_146, RQG_n, __A08_1___Q2_n, __A08_NET_144, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8028(__A08_NET_137, RL02_n_U8028_2, __A08_NET_138, __A08_1___Z2_n_U8028_4, __A08_NET_139, RL02_n_U8028_6, GND, RL02_n_U8028_8, __A08_NET_183, __A08_1___G2_n_U8028_10, __A08_NET_163, __A08_1___G2_n_U8028_12, __A08_NET_178, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8029(__A08_NET_145, WZG_n, WL02_n, __A08_NET_138, __A08_NET_145, __A08_NET_148, GND, __A08_1___Z2_n, CZG, __A08_NET_148, RZG_n, __A08_1___Z2_n, __A08_NET_147, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8030(__A08_NET_173, WBG_n, WL02_n, __A08_1___B2_n, __A08_NET_173, __A08_NET_180, GND, __A08_1___B2_n, CBG, __A08_NET_180, RBLG_n, __A08_1___B2_n, __A08_NET_181, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U8031(__A08_NET_181, __A08_NET_182, __A08_NET_177, __A08_NET_179, G02, __A08_NET_178, GND, __A08_NET_265, GND, XUY06_n, __XUY04_n, __A08_NET_183, __A08_NET_161, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8032(__A08_NET_182, __A08_NET_180, RCG_n, __A08_NET_165, WL01_n, WG3G_n, GND, WL03_n, WG4G_n, __A08_NET_164, L2GDG_n, L01_n, __A08_NET_177, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8033(__A08_NET_179, WG1G_n, WL02_n, G02, __A08_1___G2_n, CGG, GND, RGG_n, __A08_1___G2_n, __A08_NET_161, RGG_n, __G04_n, __A08_NET_255, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U8034(__A08_1___G2_n, GEM02, RL02_n, WL02, WL02, WL02_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8035(__A08_NET_297, A2XG_n, __A08_2___A1_n, __A08_NET_298, WYLOG_n, WL03_n, GND, WL02_n, WYDG_n, __A08_NET_293, __A08_2__Y1_n, CUG, __A08_2__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8036(MONEX, __A08_NET_297, __A08_2__X1_n, CLXC, CUG, __A08_2__X1, GND, __A08_2__Y1_n, __A08_NET_298, __A08_NET_293, __A08_2__Y1, __A08_2__X1_n, __A08_2__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8037(__A08_NET_302, __A08_2__X1_n, __A08_2__Y1_n, __XUY03_n, __A08_2__X1, __A08_2__Y1, GND, __A08_NET_302, __XUY03_n, __A08_NET_299, __A08_NET_302, SUMA03_n, __A08_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U8038(__A08_NET_310, __A08_NET_309, SUMA03_n, SUMB03_n, RULOG_n, __A08_NET_281, GND, __A08_NET_285, XUY05_n, __XUY03_n, __CI03_n, __A08_NET_311, G03, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U8039(__CI03_n, __A08_NET_300, __A08_2___G1_n, GEM03, RL03_n, WL03, GND, WL03_n, WL03,  ,  , __A08_NET_247, __A08_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8040(SUMB03_n, __A08_NET_299, __A08_NET_300, __A08_NET_284, WAG_n, WL03_n, GND, WL05_n, WALSG_n, __A08_NET_286, __A08_2___A1_n, CAG, __A08_NET_282, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8041(__A08_NET_285, CO06_U8041_2, __A08_NET_280, RL03_n_U8041_4, __A08_NET_289, __L03_n_U8041_6, GND, __A08_2___Z1_n_U8041_8, __A08_NET_313, RL03_n_U8041_10, __A08_NET_314, RL03_n_U8041_12, __A08_NET_315, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8042(__A08_NET_284, __A08_NET_286, __A08_NET_281, __A08_NET_279, CH03, __A08_NET_280, GND, __A08_NET_289, __A08_NET_283, __A08_NET_291, __A08_NET_292, __A08_2___A1_n, __A08_NET_282, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8043(__A08_NET_279, RAG_n, __A08_2___A1_n, __A08_NET_283, WLG_n, WL03_n, GND, G06_n, G2LSG_n, __A08_NET_291, __L03_n, CLG1G, __A08_NET_292, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8044(__A08_NET_249, __A08_2___SUMA2, __A08_2___SUMA2, __A08_2___SUMB2, RULOG_n, __A08_NET_248, GND, __A08_2___RL_OUT_1, RLG_n, __L03_n, GND, CI05_n, __CO04, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8045( ,  ,  , __A08_NET_288, WQG_n, WL03_n, GND, __A08_NET_288, __A08_NET_287, __A08_2___Q1_n, __A08_2___Q1_n, CQG, __A08_NET_287, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8046(__A08_NET_290, RQG_n, __A08_2___Q1_n, __A08_NET_316, WZG_n, WL03_n, GND, __A08_NET_316, __A08_NET_317, __A08_NET_313, __A08_2___Z1_n, CZG, __A08_NET_317, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U8047(__A08_NET_312, RZG_n, __A08_2___Z1_n, __A08_NET_322, WBG_n, WL03_n, GND, __A08_NET_322, __A08_NET_321, __A08_2___B1_n, __A08_2___B1_n, CBG, __A08_NET_321, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8048(__A08_NET_319, RBLG_n, __A08_2___B1_n, __A08_NET_318, __A08_NET_321, RCG_n, GND, WL02_n, WG3G_n, __A08_NET_307, WL04_n, WG4G_n, __A08_NET_306, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8049(__A08_2___RL_OUT_1, __A08_NET_290, MDT03, R1C, R15, __A08_NET_315, GND, __A08_NET_320, __A08_NET_319, __A08_NET_318, __A08_NET_303, __A08_NET_314, __A08_NET_312, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8050(__A08_NET_265, CO06_U8050_2, __A08_NET_320, RL03_n_U8050_4, __A08_NET_308, __A08_2___G1_n_U8050_6, GND, __A08_2___G1_n_U8050_8, __A08_NET_311, RL04_n_U8050_10, __A08_NET_235, L04_n_U8050_12, __A08_NET_236, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8051(__A08_NET_310, L2GDG_n, L02_n, __A08_NET_309, WG1G_n, WL03_n, GND, __A08_2___G1_n, CGG, G03, RGG_n, __A08_2___G1_n, __A08_NET_303, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U8052(__A08_NET_308, G03ED, SA03, __A08_NET_307, __A08_NET_306,  , GND,  , G04ED, SA04, __A08_NET_271, __A08_NET_258, __A08_NET_257, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8053(__A08_NET_250, A2XG_n, __A08_2___A2_n, __A08_NET_254, WYLOG_n, WL04_n, GND, WL03_n, WYDG_n, __A08_NET_253, __A08_2__Y2_n, CUG, __A08_2__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8054(MONEX, __A08_NET_250, __A08_2__X2_n, CLXC, CUG, __A08_2__X2, GND, __A08_2__Y2_n, __A08_NET_254, __A08_NET_253, __A08_2__Y2, __A08_2__X2_n, __A08_2__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8055(__A08_NET_249, __A08_2__X2_n, __A08_2__Y2_n, __XUY04_n, __A08_2__X2, __A08_2__Y2, GND,  ,  ,  , __A08_NET_249, __XUY04_n, __A08_NET_243, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8056(__A08_2___SUMB2, __A08_NET_243, __A08_NET_247, __A08_NET_251, WAG_n, WL04_n, GND, WL06_n, WALSG_n, __A08_NET_252, __A08_2___A2_n, CAG, __A08_NET_234, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U8057(__A08_NET_251, __A08_NET_252, __A08_NET_248, __A08_NET_233, CH04, __A08_NET_235, GND, __A08_NET_236, __A08_NET_270, __A08_NET_266, __A08_NET_269, __A08_2___A2_n, __A08_NET_234, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8058(__A08_NET_233, RAG_n, __A08_2___A2_n, __A08_NET_270, WLG_n, WL04_n, GND, G07_n, G2LSG_n, __A08_NET_266, L04_n, CLG1G, __A08_NET_269, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U8059(RLG_n, L04_n, __A08_2___RL_OUT_2, __A08_NET_237, __A08_NET_240, __A08_NET_230, GND, __A08_NET_232, MDT04, R1C, R15, __A08_2___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8060(__A08_NET_268, WQG_n, WL04_n, __A08_2___Q2_n, __A08_NET_268, __A08_NET_238, GND, __A08_2___Q2_n, CQG, __A08_NET_238, RQG_n, __A08_2___Q2_n, __A08_NET_237, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U8061(__A08_NET_230, RL04_n_U8061_2, __A08_NET_231, __A08_2___Z2_n_U8061_4, __A08_NET_232, RL04_n_U8061_6, GND, RL04_n_U8061_8, __A08_NET_278, __G04_n_U8061_10, __A08_NET_257, __G04_n_U8061_12, __A08_NET_273, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8062(__A08_NET_239, WZG_n, WL04_n, __A08_NET_231, __A08_NET_239, __A08_NET_241, GND, __A08_2___Z2_n, CZG, __A08_NET_241, RZG_n, __A08_2___Z2_n, __A08_NET_240, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U8063(__A08_NET_267, WBG_n, WL04_n, __A08_2___B2_n, __A08_NET_267, __A08_NET_275, GND, __A08_2___B2_n, CBG, __A08_NET_275, RBLG_n, __A08_2___B2_n, __A08_NET_277, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U8064(__A08_NET_276, __A08_NET_275, RCG_n, __A08_NET_271, WL03_n, WG3G_n, GND, WL05_n, WG4G_n, __A08_NET_258, L2GDG_n, __L03_n, __A08_NET_272, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U8065(__G04_n, GEM04, RL04_n, WL04, WL04, WL04_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U8066(SUMA01_n, __A08_NET_209, XUY01_n, CI01_n, GND,  , GND,  , __A08_NET_155, XUY02_n, __A08_1___CI_INTERNAL, WHOMP, SUMA02_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U8067(SUMA03_n, __A08_NET_302, __XUY03_n, __CI03_n, GND,  , GND,  , __A08_NET_249, __XUY04_n, __A08_2___CI_INTERNAL, WHOMP, __A08_2___SUMA2, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U8068(RL01_n, MWL01_U8068_2, RL02_n, MWL02_U8068_4, RL03_n, MWL03_U8068_6, GND, MWL04_U8068_8, RL04_n,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9001(__A09_NET_196, A2XG_n, __A09_1___A1_n, __A09_NET_198, WYLOG_n, WL05_n, GND, WL04_n, WYDG_n, __A09_NET_191, __A09_1__Y1_n, CUG, __A09_1__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9002(MONEX, __A09_NET_196, __A09_1__X1_n, CLXC, CUG, __A09_1__X1, GND, __A09_1__Y1_n, __A09_NET_198, __A09_NET_191, __A09_1__Y1, __A09_1__X1_n, __A09_1__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9003(__A09_NET_202, __A09_1__X1_n, __A09_1__Y1_n, XUY05_n, __A09_1__X1, __A09_1__Y1, GND, __A09_NET_202, XUY05_n, __A09_NET_200, __A09_NET_202, __A09_1___SUMA1, __A09_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9004(__A09_NET_270, __A09_NET_269, __A09_1___SUMA1, __A09_1___SUMB1, RULOG_n, __A09_NET_179, GND, __A09_NET_183, __XUY07_n, XUY05_n, CI05_n, __A09_NET_271, __A09_NET_248, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U9005(CI05_n, __A09_NET_199, G05_n, GEM05, RL05_n, WL05, GND, WL05_n, WL05,  ,  , __A09_NET_147, __A09_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9006(__A09_1___SUMB1, __A09_NET_200, __A09_NET_199, __A09_NET_182, WAG_n, WL05_n, GND, WL07_n, WALSG_n, __A09_NET_184, __A09_1___A1_n, CAG, __A09_NET_180, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9007(__A09_NET_183, __CO08_U9007_2, __A09_NET_178, RL05_n_U9007_4, __A09_NET_187, __L05_n_U9007_6, GND, __A09_1___Z1_n_U9007_8, __A09_NET_214, RL05_n_U9007_10, __A09_NET_213, RL05_n_U9007_12, __A09_NET_215, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9008(__A09_NET_177, RAG_n, __A09_1___A1_n, __A09_NET_181, WLG_n, WL05_n, GND, __G08_n, G2LSG_n, __A09_NET_189, __L05_n, CLG1G, __A09_NET_190, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9009(__A09_NET_267, WG1G_n, WL08_n, __A09_NET_186, WQG_n, WL05_n, GND, __A09_NET_186, __A09_NET_185, __A09_1___Q1_n, __A09_1___Q1_n, CQG, __A09_NET_185, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9010(__A09_NET_188, RQG_n, __A09_1___Q1_n, __A09_NET_216, WZG_n, WL05_n, GND, __A09_NET_216, __A09_NET_217, __A09_NET_214, __A09_1___Z1_n, CZG, __A09_NET_217, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9011(__A09_1___RL_OUT_1, __A09_NET_188, MDT05, R1C, GND, __A09_NET_215, GND, __A09_NET_220, __A09_NET_219, __A09_NET_218, __A09_NET_203, __A09_NET_213, __A09_NET_212, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9012(__A09_NET_212, RZG_n, __A09_1___Z1_n, __A09_NET_221, WBG_n, WL05_n, GND, __A09_NET_221, __A09_NET_222, __A09_1___B1_n, __A09_1___B1_n, CBG, __A09_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9013(__A09_NET_164, __CO08_U9013_2, __A09_NET_220, RL05_n_U9013_4, __A09_NET_208, G05_n_U9013_6, GND, G05_n_U9013_8, __A09_NET_211, RL06_n_U9013_10, __A09_NET_135, __L06_n_U9013_12, __A09_NET_136, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9014(__A09_NET_219, RBLG_n, __A09_1___B1_n, __A09_NET_218, __A09_NET_222, RCG_n, GND, WL04_n, WG3G_n, __A09_NET_207, WL06_n, WG4G_n, __A09_NET_206, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9015(__A09_NET_182, __A09_NET_184, __A09_NET_179, __A09_NET_177, CH05, __A09_NET_178, GND, __A09_NET_187, __A09_NET_181, __A09_NET_189, __A09_NET_190, __A09_1___A1_n, __A09_NET_180, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9016(__A09_NET_210, L2GDG_n, L04_n, __A09_NET_209, WG1G_n, WL05_n, GND, G05_n, CGG, G05, RGG_n, G05_n, __A09_NET_203, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U9017(__A09_NET_210, __A09_NET_209, GND, __XUY08_n, XUY06_n, __A09_NET_164, GND, __A09_1___RL_OUT_1, RLG_n, __L05_n, GND, __A09_NET_211, G05, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U9018(__A09_NET_208, G05ED, SA05, __A09_NET_207, __A09_NET_206,  , GND,  , G06ED, SA06, __A09_NET_158, __A09_NET_157, __A09_NET_156, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9019(__A09_NET_149, A2XG_n, __A09_1___A2_n, __A09_NET_153, WYLOG_n, WL06_n, GND, WL05_n, WYDG_n, __A09_NET_152, __A09_1__Y2_n, CUG, __A09_1__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9020(MONEX, __A09_NET_149, __A09_1__X2_n, CLXC, CUG, __A09_1__X2, GND, __A09_1__Y2_n, __A09_NET_153, __A09_NET_152, __A09_1__Y2, __A09_1__X2_n, __A09_1__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9021(__A09_NET_148, __A09_1__X2_n, __A09_1__Y2_n, XUY06_n, __A09_1__X2, __A09_1__Y2, GND, __G08_n, CGG, G08, __A09_NET_148, XUY06_n, __A09_NET_143, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U9022(__A09_NET_265, __A09_NET_267, __A09_NET_148, __A09_1___SUMA2, CO06, __CI07_n, GND, __A09_NET_197, __A09_1___SUMA2, __A09_1___SUMB2, RULOG_n, __A09_NET_266, G08, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9023(__A09_1___SUMB2, __A09_NET_143, __A09_NET_147, __A09_NET_150, WAG_n, WL06_n, GND, WL08_n, WALSG_n, __A09_NET_151, __A09_1___A2_n, CAG, __A09_NET_134, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9024(__A09_NET_150, __A09_NET_151, __A09_NET_197, __A09_NET_133, CH06, __A09_NET_135, GND, __A09_NET_136, __A09_NET_168, __A09_NET_165, __A09_NET_169, __A09_1___A2_n, __A09_NET_134, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9025(__A09_NET_133, RAG_n, __A09_1___A2_n, __A09_NET_168, WLG_n, WL06_n, GND, G09_n, G2LSG_n, __A09_NET_165, __L06_n, CLG1G, __A09_NET_169, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9026(RLG_n, __L06_n, __A09_1___RL_OUT_2, __A09_NET_137, __A09_NET_140, __A09_NET_130, GND, __A09_NET_132, MDT06, R1C, GND, __A09_1___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9027(__A09_NET_167, WQG_n, WL06_n, __A09_1___Q2_n, __A09_NET_167, __A09_NET_139, GND, __A09_1___Q2_n, CQG, __A09_NET_139, RQG_n, __A09_1___Q2_n, __A09_NET_137, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9028(__A09_NET_130, RL06_n_U9028_2, __A09_NET_131, __A09_1___Z2_n_U9028_4, __A09_NET_132, RL06_n_U9028_6, GND, RL06_n_U9028_8, __A09_NET_176, G06_n_U9028_10, __A09_NET_156, G06_n_U9028_12, __A09_NET_171, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9029(__A09_NET_138, WZG_n, WL06_n, __A09_NET_131, __A09_NET_138, __A09_NET_141, GND, __A09_1___Z2_n, CZG, __A09_NET_141, RZG_n, __A09_1___Z2_n, __A09_NET_140, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9030(__A09_NET_166, WBG_n, WL06_n, __A09_1___B2_n, __A09_NET_166, __A09_NET_173, GND, __A09_1___B2_n, CBG, __A09_NET_173, RBLG_n, __A09_1___B2_n, __A09_NET_174, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U9031(__A09_NET_174, __A09_NET_175, __A09_NET_170, __A09_NET_172, G06, __A09_NET_171, GND, __A09_NET_258, GND, XUY10_n, __XUY08_n, __A09_NET_176, __A09_NET_154, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9032(__A09_NET_175, __A09_NET_173, RCG_n, __A09_NET_158, WL05_n, WG3G_n, GND, WL07_n, WG4G_n, __A09_NET_157, L2GDG_n, __L05_n, __A09_NET_170, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9033(__A09_NET_172, WG1G_n, WL06_n, G06, G06_n, CGG, GND, RGG_n, G06_n, __A09_NET_154, RGG_n, __G08_n, __A09_NET_248, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U9034(G06_n, GEM06, RL06_n, WL06, WL06, WL06_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9035(__A09_NET_290, A2XG_n, __A09_2___A1_n, __A09_NET_291, WYLOG_n, WL07_n, GND, WL06_n, WYDG_n, __A09_NET_286, __A09_2__Y1_n, CUG, __A09_2__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9036(MONEX, __A09_NET_290, __A09_2__X1_n, CLXC, CUG, __A09_2__X1, GND, __A09_2__Y1_n, __A09_NET_291, __A09_NET_286, __A09_2__Y1, __A09_2__X1_n, __A09_2__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9037(__A09_NET_295, __A09_2__X1_n, __A09_2__Y1_n, __XUY07_n, __A09_2__X1, __A09_2__Y1, GND, __A09_NET_295, __XUY07_n, __A09_NET_292, __A09_NET_295, __A09_2___SUMA1, __A09_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U9038(__A09_NET_303, __A09_NET_302, __A09_2___SUMA1, __A09_2___SUMB1, RULOG_n, __A09_NET_274, GND, __A09_NET_278, XUY09_n, __XUY07_n, __CI07_n, __A09_NET_304, G07, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U9039(__CI07_n, __A09_NET_293, G07_n, GEM07, __A09_2___RL1_n, WL07, GND, WL07_n, WL07,  ,  , __A09_NET_240, __A09_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9040(__A09_2___SUMB1, __A09_NET_292, __A09_NET_293, __A09_NET_277, WAG_n, WL07_n, GND, WL09_n, WALSG_n, __A09_NET_279, __A09_2___A1_n, CAG, __A09_NET_275, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9041(__A09_NET_278, CO10_U9041_2, __A09_NET_273, __A09_2___RL1_n_U9041_4, __A09_NET_282, __L07_n_U9041_6, GND, __A09_2___Z1_n_U9041_8, __A09_NET_306, __A09_2___RL1_n_U9041_10, __A09_NET_307, __A09_2___RL1_n_U9041_12, __A09_NET_308, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9042(__A09_NET_277, __A09_NET_279, __A09_NET_274, __A09_NET_272, CH07, __A09_NET_273, GND, __A09_NET_282, __A09_NET_276, __A09_NET_284, __A09_NET_285, __A09_2___A1_n, __A09_NET_275, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9043(__A09_NET_272, RAG_n, __A09_2___A1_n, __A09_NET_276, WLG_n, WL07_n, GND, G10_n, G2LSG_n, __A09_NET_284, __L07_n, CLG1G, __A09_NET_285, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9044(__A09_NET_242, __A09_2___SUMA2, __A09_2___SUMA2, __A09_2___SUMB2, RULOG_n, __A09_NET_241, GND, __A09_2___RL_OUT_1, RLG_n, __L07_n, GND, CI09_n, __CO08, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9045( ,  ,  , __A09_NET_281, WQG_n, WL07_n, GND, __A09_NET_281, __A09_NET_280, __A09_2___Q1_n, __A09_2___Q1_n, CQG, __A09_NET_280, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9046(__A09_NET_283, RQG_n, __A09_2___Q1_n, __A09_NET_309, WZG_n, WL07_n, GND, __A09_NET_309, __A09_NET_310, __A09_NET_306, __A09_2___Z1_n, CZG, __A09_NET_310, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U9047(__A09_NET_305, RZG_n, __A09_2___Z1_n, __A09_NET_315, WBG_n, WL07_n, GND, __A09_NET_315, __A09_NET_314, __A09_2___B1_n, __A09_2___B1_n, CBG, __A09_NET_314, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9048(__A09_NET_312, RBLG_n, __A09_2___B1_n, __A09_NET_311, __A09_NET_314, RCG_n, GND, WL06_n, WG3G_n, __A09_NET_300, WL08_n, WG4G_n, __A09_NET_299, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9049(__A09_2___RL_OUT_1, __A09_NET_283, MDT07, R1C, GND, __A09_NET_308, GND, __A09_NET_313, __A09_NET_312, __A09_NET_311, __A09_NET_296, __A09_NET_307, __A09_NET_305, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9050(__A09_NET_258, CO10_U9050_2, __A09_NET_313, __A09_2___RL1_n_U9050_4, __A09_NET_301, G07_n_U9050_6, GND, G07_n_U9050_8, __A09_NET_304, __A09_2___RL2_n_U9050_10, __A09_NET_228, L08_n_U9050_12, __A09_NET_229, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9051(__A09_NET_303, L2GDG_n, __L06_n, __A09_NET_302, WG1G_n, WL07_n, GND, G07_n, CGG, G07, RGG_n, G07_n, __A09_NET_296, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U9052(__A09_NET_301, G07ED, SA07, __A09_NET_300, __A09_NET_299,  , GND,  , GND, SA08, __A09_NET_264, __A09_NET_251, __A09_NET_250, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9053(__A09_NET_243, A2XG_n, __A09_2___A2_n, __A09_NET_247, WYLOG_n, WL08_n, GND, WL07_n, WYDG_n, __A09_NET_246, __A09_2__Y2_n, CUG, __A09_2__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9054(MONEX, __A09_NET_243, __A09_2__X2_n, CLXC, CUG, __A09_2__X2, GND, __A09_2__Y2_n, __A09_NET_247, __A09_NET_246, __A09_2__Y2, __A09_2__X2_n, __A09_2__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9055(__A09_NET_242, __A09_2__X2_n, __A09_2__Y2_n, __XUY08_n, __A09_2__X2, __A09_2__Y2, GND,  ,  ,  , __A09_NET_242, __XUY08_n, __A09_NET_236, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9056(__A09_2___SUMB2, __A09_NET_236, __A09_NET_240, __A09_NET_244, WAG_n, WL08_n, GND, WL10_n, WALSG_n, __A09_NET_245, __A09_2___A2_n, CAG, __A09_NET_227, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U9057(__A09_NET_244, __A09_NET_245, __A09_NET_241, __A09_NET_226, CH08, __A09_NET_228, GND, __A09_NET_229, __A09_NET_263, __A09_NET_259, __A09_NET_262, __A09_2___A2_n, __A09_NET_227, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9058(__A09_NET_226, RAG_n, __A09_2___A2_n, __A09_NET_263, WLG_n, WL08_n, GND, G11_n, G2LSG_n, __A09_NET_259, L08_n, CLG1G, __A09_NET_262, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U9059(RLG_n, L08_n, __A09_2___RL_OUT_2, __A09_NET_230, __A09_NET_233, __A09_NET_223, GND, __A09_NET_225, MDT08, R1C, GND, __A09_2___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9060(__A09_NET_261, WQG_n, WL08_n, __A09_2___Q2_n, __A09_NET_261, __A09_NET_231, GND, __A09_2___Q2_n, CQG, __A09_NET_231, RQG_n, __A09_2___Q2_n, __A09_NET_230, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U9061(__A09_NET_223, __A09_2___RL2_n_U9061_2, __A09_NET_224, __A09_2___Z2_n_U9061_4, __A09_NET_225, __A09_2___RL2_n_U9061_6, GND, __A09_2___RL2_n_U9061_8, __A09_NET_271, __G08_n_U9061_10, __A09_NET_250, __G08_n_U9061_12, __A09_NET_266, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9062(__A09_NET_232, WZG_n, WL08_n, __A09_NET_224, __A09_NET_232, __A09_NET_234, GND, __A09_2___Z2_n, CZG, __A09_NET_234, RZG_n, __A09_2___Z2_n, __A09_NET_233, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U9063(__A09_NET_260, WBG_n, WL08_n, __A09_2___B2_n, __A09_NET_260, __A09_NET_268, GND, __A09_2___B2_n, CBG, __A09_NET_268, RBLG_n, __A09_2___B2_n, __A09_NET_270, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U9064(__A09_NET_269, __A09_NET_268, RCG_n, __A09_NET_264, WL07_n, WG3G_n, GND, WL09_n, WG4G_n, __A09_NET_251, L2GDG_n, __L07_n, __A09_NET_265, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U9065(__G08_n, GEM08, __A09_2___RL2_n, WL08, WL08, WL08_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U9066(__A09_1___SUMA1, __A09_NET_202, XUY05_n, CI05_n, GND,  , GND,  , __A09_NET_148, XUY06_n, __A09_1___CI_INTERNAL, GND, __A09_1___SUMA2, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U9067(__A09_2___SUMA1, __A09_NET_295, __XUY07_n, __CI07_n, WHOMP,  , GND,  , __A09_NET_242, __XUY08_n, __A09_2___CI_INTERNAL, GND, __A09_2___SUMA2, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U9068(RL05_n, MWL05_U9068_2, RL06_n, MWL06_U9068_4, __A09_2___RL1_n, MWL07_U9068_6, GND, MWL08_U9068_8, __A09_2___RL2_n,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10001(__A10_NET_195, A2XG_n, __A10_1___A1_n, __A10_NET_197, WYLOG_n, WL09_n, GND, WL08_n, WYDG_n, __A10_NET_190, __A10_1__Y1_n, CUG, __A10_1__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10002(MONEX, __A10_NET_195, __A10_1__X1_n, CLXC, CUG, __A10_1__X1, GND, __A10_1__Y1_n, __A10_NET_197, __A10_NET_190, __A10_1__Y1, __A10_1__X1_n, __A10_1__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10003(__A10_NET_201, __A10_1__X1_n, __A10_1__Y1_n, XUY09_n, __A10_1__X1, __A10_1__Y1, GND, __A10_NET_201, XUY09_n, __A10_NET_199, __A10_NET_201, __A10_1___SUMA1, __A10_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U10004(__A10_NET_269, __A10_NET_268, __A10_1___SUMA1, __A10_1___SUMB1, RULOG_n, __A10_NET_178, GND, __A10_NET_182, __XUY11_n, XUY09_n, CI09_n, __A10_NET_270, __A10_NET_247, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U10005(CI09_n, __A10_NET_198, G09_n, GEM09, RL09_n, WL09, GND, WL09_n, WL09,  ,  , __A10_NET_146, __A10_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10006(__A10_1___SUMB1, __A10_NET_199, __A10_NET_198, __A10_NET_181, WAG_n, WL09_n, GND, WL11_n, WALSG_n, __A10_NET_183, __A10_1___A1_n, CAG, __A10_NET_179, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U10007(__A10_NET_182, __CO12_U10007_2, __A10_NET_177, RL09_n_U10007_4, __A10_NET_186, __L09_n_U10007_6, GND, __A10_1___Z1_n_U10007_8, __A10_NET_213, RL09_n_U10007_10, __A10_NET_212, RL09_n_U10007_12, __A10_NET_214, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10008(__A10_NET_176, RAG_n, __A10_1___A1_n, __A10_NET_180, WLG_n, WL09_n, GND, __G12_n, G2LSG_n, __A10_NET_188, __L09_n, CLG1G, __A10_NET_189, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10009(__A10_NET_266, WG1G_n, WL12_n, __A10_NET_185, WQG_n, WL09_n, GND, __A10_NET_185, __A10_NET_184, __A10_1___Q1_n, __A10_1___Q1_n, CQG, __A10_NET_184, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10010(__A10_NET_187, RQG_n, __A10_1___Q1_n, __A10_NET_215, WZG_n, WL09_n, GND, __A10_NET_215, __A10_NET_216, __A10_NET_213, __A10_1___Z1_n, CZG, __A10_NET_216, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U10011(__A10_1___RL_OUT_1, __A10_NET_187, MDT09, R1C, GND, __A10_NET_214, GND, __A10_NET_219, __A10_NET_218, __A10_NET_217, __A10_NET_202, __A10_NET_212, __A10_NET_211, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10012(__A10_NET_211, RZG_n, __A10_1___Z1_n, __A10_NET_220, WBG_n, WL09_n, GND, __A10_NET_220, __A10_NET_221, __A10_1___B1_n, __A10_1___B1_n, CBG, __A10_NET_221, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U10013(__A10_NET_163, __CO12_U10013_2, __A10_NET_219, RL09_n_U10013_4, __A10_NET_207, G09_n_U10013_6, GND, G09_n_U10013_8, __A10_NET_210, RL10_n_U10013_10, __A10_NET_134, __L10_n_U10013_12, __A10_NET_135, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10014(__A10_NET_218, RBLG_n, __A10_1___B1_n, __A10_NET_217, __A10_NET_221, RCG_n, GND, WL08_n, WG3G_n, __A10_NET_206, WL10_n, WG4G_n, __A10_NET_205, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10015(__A10_NET_181, __A10_NET_183, __A10_NET_178, __A10_NET_176, CH09, __A10_NET_177, GND, __A10_NET_186, __A10_NET_180, __A10_NET_188, __A10_NET_189, __A10_1___A1_n, __A10_NET_179, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10016(__A10_NET_209, L2GDG_n, L08_n, __A10_NET_208, WG1G_n, WL09_n, GND, G09_n, CGG, G09, RGG_n, G09_n, __A10_NET_202, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U10017(__A10_NET_209, __A10_NET_208, WHOMPA, __XUY12_n, XUY10_n, __A10_NET_163, GND, __A10_1___RL_OUT_1, RLG_n, __L09_n, GND, __A10_NET_210, G09, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U10018(__A10_NET_207, GND, SA09, __A10_NET_206, __A10_NET_205,  , GND,  , GND, SA10, __A10_NET_157, __A10_NET_156, __A10_NET_155, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10019(__A10_NET_148, A2XG_n, __A10_1___A2_n, __A10_NET_152, WYLOG_n, WL10_n, GND, WL09_n, WYDG_n, __A10_NET_151, __A10_1__Y2_n, CUG, __A10_1__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10020(MONEX, __A10_NET_148, __A10_1__X2_n, CLXC, CUG, __A10_1__X2, GND, __A10_1__Y2_n, __A10_NET_152, __A10_NET_151, __A10_1__Y2, __A10_1__X2_n, __A10_1__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10021(__A10_NET_147, __A10_1__X2_n, __A10_1__Y2_n, XUY10_n, __A10_1__X2, __A10_1__Y2, GND, __G12_n, CGG, G12, __A10_NET_147, XUY10_n, __A10_NET_142, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U10022(__A10_NET_264, __A10_NET_266, __A10_NET_147, __A10_1___SUMA2, CO10, __CI11_n, GND, __A10_NET_196, __A10_1___SUMA2, __A10_1___SUMB2, RULOG_n, __A10_NET_265, G12, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10023(__A10_1___SUMB2, __A10_NET_142, __A10_NET_146, __A10_NET_149, WAG_n, WL10_n, GND, WL12_n, WALSG_n, __A10_NET_150, __A10_1___A2_n, CAG, __A10_NET_133, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10024(__A10_NET_149, __A10_NET_150, __A10_NET_196, __A10_NET_132, CH10, __A10_NET_134, GND, __A10_NET_135, __A10_NET_167, __A10_NET_164, __A10_NET_168, __A10_1___A2_n, __A10_NET_133, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10025(__A10_NET_132, RAG_n, __A10_1___A2_n, __A10_NET_167, WLG_n, WL10_n, GND, G13_n, G2LSG_n, __A10_NET_164, __L10_n, CLG1G, __A10_NET_168, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U10026(RLG_n, __L10_n, __A10_1___RL_OUT_2, __A10_NET_136, __A10_NET_139, __A10_NET_129, GND, __A10_NET_131, MDT10, R1C, GND, __A10_1___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10027(__A10_NET_166, WQG_n, WL10_n, __A10_1___Q2_n, __A10_NET_166, __A10_NET_138, GND, __A10_1___Q2_n, CQG, __A10_NET_138, RQG_n, __A10_1___Q2_n, __A10_NET_136, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U10028(__A10_NET_129, RL10_n_U10028_2, __A10_NET_130, __A10_1___Z2_n_U10028_4, __A10_NET_131, RL10_n_U10028_6, GND, RL10_n_U10028_8, __A10_NET_175, G10_n_U10028_10, __A10_NET_155, G10_n_U10028_12, __A10_NET_170, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10029(__A10_NET_137, WZG_n, WL10_n, __A10_NET_130, __A10_NET_137, __A10_NET_140, GND, __A10_1___Z2_n, CZG, __A10_NET_140, RZG_n, __A10_1___Z2_n, __A10_NET_139, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10030(__A10_NET_165, WBG_n, WL10_n, __A10_1___B2_n, __A10_NET_165, __A10_NET_172, GND, __A10_1___B2_n, CBG, __A10_NET_172, RBLG_n, __A10_1___B2_n, __A10_NET_173, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U10031(__A10_NET_173, __A10_NET_174, __A10_NET_169, __A10_NET_171, G10, __A10_NET_170, GND, __A10_NET_257, GND, XUY14_n, __XUY12_n, __A10_NET_175, __A10_NET_153, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10032(__A10_NET_174, __A10_NET_172, RCG_n, __A10_NET_157, WL09_n, WG3G_n, GND, WL11_n, WG4G_n, __A10_NET_156, L2GDG_n, __L09_n, __A10_NET_169, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10033(__A10_NET_171, WG1G_n, WL10_n, G10, G10_n, CGG, GND, RGG_n, G10_n, __A10_NET_153, RGG_n, __G12_n, __A10_NET_247, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U10034(G10_n, GEM10, RL10_n, WL10, WL10, WL10_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10035(__A10_NET_289, A2XG_n, __A10_2___A1_n, __A10_NET_290, WYLOG_n, WL11_n, GND, WL10_n, WYDG_n, __A10_NET_285, __A10_2__Y1_n, CUG, __A10_2__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10036(MONEX, __A10_NET_289, __A10_2__X1_n, CLXC, CUG, __A10_2__X1, GND, __A10_2__Y1_n, __A10_NET_290, __A10_NET_285, __A10_2__Y1, __A10_2__X1_n, __A10_2__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10037(__A10_NET_294, __A10_2__X1_n, __A10_2__Y1_n, __XUY11_n, __A10_2__X1, __A10_2__Y1, GND, __A10_NET_294, __XUY11_n, __A10_NET_291, __A10_NET_294, SUMA11_n, __A10_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U10038(__A10_NET_302, __A10_NET_301, SUMA11_n, SUMB11_n, RULOG_n, __A10_NET_273, GND, __A10_NET_277, XUY13_n, __XUY11_n, __CI11_n, __A10_NET_303, G11, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U10039(__CI11_n, __A10_NET_292, G11_n, GEM11, RL11_n, WL11, GND, WL11_n, WL11,  ,  , __A10_NET_239, __A10_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10040(SUMB11_n, __A10_NET_291, __A10_NET_292, __A10_NET_276, WAG_n, WL11_n, GND, WL13_n, WALSG_n, __A10_NET_278, __A10_2___A1_n, CAG, __A10_NET_274, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U10041(__A10_NET_277, CO14_U10041_2, __A10_NET_272, RL11_n_U10041_4, __A10_NET_281, __L11_n_U10041_6, GND, __A10_2___Z1_n_U10041_8, __A10_NET_305, RL11_n_U10041_10, __A10_NET_306, RL11_n_U10041_12, __A10_NET_307, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10042(__A10_NET_276, __A10_NET_278, __A10_NET_273, __A10_NET_271, CH11, __A10_NET_272, GND, __A10_NET_281, __A10_NET_275, __A10_NET_283, __A10_NET_284, __A10_2___A1_n, __A10_NET_274, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10043(__A10_NET_271, RAG_n, __A10_2___A1_n, __A10_NET_275, WLG_n, WL11_n, GND, G14_n, G2LSG_n, __A10_NET_283, __L11_n, CLG1G, __A10_NET_284, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U10044(__A10_NET_241, SUMA12_n, SUMA12_n, SUMB12_n, RULOG_n, __A10_NET_240, GND, __A10_2___RL_OUT_1, RLG_n, __L11_n, GND, CI13_n, __CO12, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10045( ,  ,  , __A10_NET_280, WQG_n, WL11_n, GND, __A10_NET_280, __A10_NET_279, __A10_2___Q1_n, __A10_2___Q1_n, CQG, __A10_NET_279, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10046(__A10_NET_282, RQG_n, __A10_2___Q1_n, __A10_NET_308, WZG_n, WL11_n, GND, __A10_NET_308, __A10_NET_309, __A10_NET_305, __A10_2___Z1_n, CZG, __A10_NET_309, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U10047(__A10_NET_304, RZG_n, __A10_2___Z1_n, __A10_NET_314, WBG_n, WL11_n, GND, __A10_NET_314, __A10_NET_313, __A10_2___B1_n, __A10_2___B1_n, CBG, __A10_NET_313, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10048(__A10_NET_311, RBHG_n, __A10_2___B1_n, __A10_NET_310, __A10_NET_313, RCG_n, GND, WL10_n, WG3G_n, __A10_NET_299, WL12_n, WG4G_n, __A10_NET_298, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U10049(__A10_2___RL_OUT_1, __A10_NET_282, MDT11, R1C, GND, __A10_NET_307, GND, __A10_NET_312, __A10_NET_311, __A10_NET_310, __A10_NET_295, __A10_NET_306, __A10_NET_304, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U10050(__A10_NET_257, CO14_U10050_2, __A10_NET_312, RL11_n_U10050_4, __A10_NET_300, G11_n_U10050_6, GND, G11_n_U10050_8, __A10_NET_303, RL12_n_U10050_10, __A10_NET_227, L12_n_U10050_12, __A10_NET_228, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10051(__A10_NET_302, L2GDG_n, __L10_n, __A10_NET_301, WG1G_n, WL11_n, GND, G11_n, CGG, G11, RGG_n, G11_n, __A10_NET_295, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U10052(__A10_NET_300, GND, SA11, __A10_NET_299, __A10_NET_298,  , GND,  , GND, SA12, __A10_NET_263, __A10_NET_250, __A10_NET_249, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10053(__A10_NET_242, A2XG_n, __A10_2___A2_n, __A10_NET_246, WYLOG_n, WL12_n, GND, WL11_n, WYDG_n, __A10_NET_245, __A10_2__Y2_n, CUG, __A10_2__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10054(MONEX, __A10_NET_242, __A10_2__X2_n, CLXC, CUG, __A10_2__X2, GND, __A10_2__Y2_n, __A10_NET_246, __A10_NET_245, __A10_2__Y2, __A10_2__X2_n, __A10_2__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10055(__A10_NET_241, __A10_2__X2_n, __A10_2__Y2_n, __XUY12_n, __A10_2__X2, __A10_2__Y2, GND,  ,  ,  , __A10_NET_241, __XUY12_n, __A10_NET_235, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10056(SUMB12_n, __A10_NET_235, __A10_NET_239, __A10_NET_243, WAG_n, WL12_n, GND, WL14_n, WALSG_n, __A10_NET_244, __A10_2___A2_n, CAG, __A10_NET_226, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U10057(__A10_NET_243, __A10_NET_244, __A10_NET_240, __A10_NET_225, CH12, __A10_NET_227, GND, __A10_NET_228, __A10_NET_262, __A10_NET_258, __A10_NET_261, __A10_2___A2_n, __A10_NET_226, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10058(__A10_NET_225, RAG_n, __A10_2___A2_n, __A10_NET_262, WLG_n, WL12_n, GND, G15_n, G2LSG_n, __A10_NET_258, L12_n, CLG1G, __A10_NET_261, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U10059(RLG_n, L12_n, __A10_2___RL_OUT_2, __A10_NET_229, __A10_NET_232, __A10_NET_222, GND, __A10_NET_224, MDT12, R1C, GND, __A10_2___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10060(__A10_NET_260, WQG_n, WL12_n, __A10_2___Q2_n, __A10_NET_260, __A10_NET_230, GND, __A10_2___Q2_n, CQG, __A10_NET_230, RQG_n, __A10_2___Q2_n, __A10_NET_229, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U10061(__A10_NET_222, RL12_n_U10061_2, __A10_NET_223, __A10_2___Z2_n_U10061_4, __A10_NET_224, RL12_n_U10061_6, GND, RL12_n_U10061_8, __A10_NET_270, __G12_n_U10061_10, __A10_NET_249, __G12_n_U10061_12, __A10_NET_265, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10062(__A10_NET_231, WZG_n, WL12_n, __A10_NET_223, __A10_NET_231, __A10_NET_233, GND, __A10_2___Z2_n, CZG, __A10_NET_233, RZG_n, __A10_2___Z2_n, __A10_NET_232, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U10063(__A10_NET_259, WBG_n, WL12_n, __A10_2___B2_n, __A10_NET_259, __A10_NET_267, GND, __A10_2___B2_n, CBG, __A10_NET_267, RBHG_n, __A10_2___B2_n, __A10_NET_269, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U10064(__A10_NET_268, __A10_NET_267, RCG_n, __A10_NET_263, WL11_n, WG3G_n, GND, WL13_n, WG4G_n, __A10_NET_250, L2GDG_n, __L11_n, __A10_NET_264, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U10065(__G12_n, GEM12, RL12_n, WL12, WL12, WL12_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U10066(__A10_1___SUMA1, __A10_NET_201, XUY09_n, CI09_n, GND,  , GND,  , __A10_NET_147, XUY10_n, __A10_1___CI_INTERNAL, GND, __A10_1___SUMA2, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U10067(SUMA11_n, __A10_NET_294, __XUY11_n, __CI11_n, GND,  , GND,  , __A10_NET_241, __XUY12_n, __A10_2___CI_INTERNAL, WHOMP, SUMA12_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U10068(RL09_n, MWL09_U10068_2, RL10_n, MWL10_U10068_4, RL11_n, MWL11_U10068_6, GND, MWL12_U10068_8, RL12_n,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11001(__A11_NET_196, A2XG_n, __A11_1___A1_n, __A11_NET_198, WYHIG_n, WL13_n, GND, WL12_n, WYDG_n, __A11_NET_191, __A11_1__Y1_n, CUG, __A11_1__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11002(MONEX, __A11_NET_196, __A11_1__X1_n, CLXC, CUG, __A11_1__X1, GND, __A11_1__Y1_n, __A11_NET_198, __A11_NET_191, __A11_1__Y1, __A11_1__X1_n, __A11_1__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11003(__A11_NET_202, __A11_1__X1_n, __A11_1__Y1_n, XUY13_n, __A11_1__X1, __A11_1__Y1, GND, __A11_NET_202, XUY13_n, __A11_NET_200, __A11_NET_202, SUMA13_n, __A11_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11004(__A11_NET_270, __A11_NET_269, SUMA13_n, SUMB13_n, RULOG_n, __A11_NET_179, GND, __A11_NET_183, __XUY15_n, XUY13_n, CI13_n, __A11_NET_271, __A11_NET_248, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11005(CI13_n, __A11_NET_199, G13_n, GEM13, RL13_n, WL13, GND, WL13_n, WL13,  ,  , __A11_NET_147, __A11_1___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11006(SUMB13_n, __A11_NET_200, __A11_NET_199, __A11_NET_182, WAG_n, WL13_n, GND, WL15_n, WALSG_n, __A11_NET_184, __A11_1___A1_n, CAG, __A11_NET_180, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11007(__A11_NET_183, __CO16_U11007_2, __A11_NET_178, RL13_n_U11007_4, __A11_NET_187, __L13_n_U11007_6, GND, __A11_1___Z1_n_U11007_8, __A11_NET_214, RL13_n_U11007_10, __A11_NET_213, RL13_n_U11007_12, __A11_NET_215, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11008(__A11_NET_177, RAG_n, __A11_1___A1_n, __A11_NET_181, WLG_n, WL13_n, GND, WL01_n, WALSG_n, __A11_NET_189, __L13_n, CLG2G, __A11_NET_190, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11009(__A11_NET_267, WG2G_n, WL16_n, __A11_NET_186, WQG_n, WL13_n, GND, __A11_NET_186, __A11_NET_185, __A11_1___Q1_n, __A11_1___Q1_n, CQG, __A11_NET_185, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11010(__A11_NET_188, RQG_n, __A11_1___Q1_n, __A11_NET_216, WZG_n, WL13_n, GND, __A11_NET_216, __A11_NET_217, __A11_NET_214, __A11_1___Z1_n, CZG, __A11_NET_217, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11011(__A11_1___RL_OUT_1, __A11_NET_188, MDT13, R1C, GND, __A11_NET_215, GND, __A11_NET_220, __A11_NET_219, __A11_NET_218, __A11_NET_203, __A11_NET_213, __A11_NET_212, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11012(__A11_NET_212, RZG_n, __A11_1___Z1_n, __A11_NET_221, WBG_n, WL13_n, GND, __A11_NET_221, __A11_NET_222, __A11_1___B1_n, __A11_1___B1_n, CBG, __A11_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11013(__A11_NET_164, __CO16_U11013_2, __A11_NET_220, RL13_n_U11013_4, __A11_NET_208, G13_n_U11013_6, GND, G13_n_U11013_8, __A11_NET_211, RL14_n_U11013_10, __A11_NET_135, __L14_n_U11013_12, __A11_NET_136, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11014(__A11_NET_219, RBHG_n, __A11_1___B1_n, __A11_NET_218, __A11_NET_222, RCG_n, GND, WL12_n, WG3G_n, __A11_NET_207, WL14_n, WG4G_n, __A11_NET_206, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11015(__A11_NET_182, __A11_NET_184, __A11_NET_179, __A11_NET_177, CH13, __A11_NET_178, GND, __A11_NET_187, __A11_NET_181, __A11_NET_189, __A11_NET_190, __A11_1___A1_n, __A11_NET_180, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11016(__A11_NET_210, L2GDG_n, L12_n, __A11_NET_209, WG1G_n, WL13_n, GND, G13_n, CGG, G13, RGG_n, G13_n, __A11_NET_203, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U11017(__A11_NET_210, __A11_NET_209, GND, __XUY16_n, XUY14_n, __A11_NET_164, GND, __A11_1___RL_OUT_1, RLG_n, __L13_n, GND, __A11_NET_211, G13, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U11018(__A11_NET_208, GND, SA13, __A11_NET_207, __A11_NET_206,  , GND,  , GND, SA14, __A11_NET_158, __A11_NET_157, __A11_NET_156, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11019(__A11_NET_149, A2XG_n, __A11_1___A2_n, __A11_NET_153, WYHIG_n, WL14_n, GND, WL13_n, WYDG_n, __A11_NET_152, __A11_1__Y2_n, CUG, __A11_1__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11020(MONEX, __A11_NET_149, __A11_1__X2_n, CLXC, CUG, __A11_1__X2, GND, __A11_1__Y2_n, __A11_NET_153, __A11_NET_152, __A11_1__Y2, __A11_1__X2_n, __A11_1__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11021(__A11_NET_148, __A11_1__X2_n, __A11_1__Y2_n, XUY14_n, __A11_1__X2, __A11_1__Y2, GND, __G16_n, CGG, G16, __A11_NET_148, XUY14_n, __A11_NET_143, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U11022(__A11_NET_265, __A11_NET_267, __A11_NET_148, SUMA14_n, CO14, __CI15_n, GND, __A11_NET_197, SUMA14_n, SUMB14_n, RULOG_n, __A11_NET_266, G16, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11023(SUMB14_n, __A11_NET_143, __A11_NET_147, __A11_NET_150, WAG_n, WL14_n, GND, WL16_n, WALSG_n, __A11_NET_151, __A11_1___A2_n, CAG, __A11_NET_134, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11024(__A11_NET_150, __A11_NET_151, __A11_NET_197, __A11_NET_133, CH14, __A11_NET_135, GND, __A11_NET_136, __A11_NET_168, __A11_NET_165, __A11_NET_169, __A11_1___A2_n, __A11_NET_134, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11025(__A11_NET_133, RAG_n, __A11_1___A2_n, __A11_NET_168, WLG_n, WL14_n, GND, WL02_n, WALSG_n, __A11_NET_165, __L14_n, CLG2G, __A11_NET_169, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11026(RLG_n, __L14_n, __A11_1___RL_OUT_2, __A11_NET_137, __A11_NET_140, __A11_NET_130, GND, __A11_NET_132, MDT14, R1C, GND, __A11_1___RL_OUT_2, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11027(__A11_NET_167, WQG_n, WL14_n, __A11_1___Q2_n, __A11_NET_167, __A11_NET_139, GND, __A11_1___Q2_n, CQG, __A11_NET_139, RQG_n, __A11_1___Q2_n, __A11_NET_137, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11028(__A11_NET_130, RL14_n_U11028_2, __A11_NET_131, __A11_1___Z2_n_U11028_4, __A11_NET_132, RL14_n_U11028_6, GND, RL14_n_U11028_8, __A11_NET_176, G14_n_U11028_10, __A11_NET_156, G14_n_U11028_12, __A11_NET_171, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11029(__A11_NET_138, WZG_n, WL14_n, __A11_NET_131, __A11_NET_138, __A11_NET_141, GND, __A11_1___Z2_n, CZG, __A11_NET_141, RZG_n, __A11_1___Z2_n, __A11_NET_140, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11030(__A11_NET_166, WBG_n, WL14_n, __A11_1___B2_n, __A11_NET_166, __A11_NET_173, GND, __A11_1___B2_n, CBG, __A11_NET_173, RBHG_n, __A11_1___B2_n, __A11_NET_174, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U11031(__A11_NET_174, __A11_NET_175, __A11_NET_170, __A11_NET_172, G14, __A11_NET_171, GND, __A11_NET_258, GND, XUY02_n, __XUY16_n, __A11_NET_176, __A11_NET_154, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11032(__A11_NET_175, __A11_NET_173, RCG_n, __A11_NET_158, WL13_n, WG3G_n, GND, WL16_n, WG4G_n, __A11_NET_157, L2GDG_n, __L13_n, __A11_NET_170, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11033(__A11_NET_172, WG1G_n, WL14_n, G14, G14_n, CGG, GND, RGG_n, G14_n, __A11_NET_154, RGG_n, __G16_n, __A11_NET_248, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11034(G14_n, GEM14, RL14_n, WL14, WL14, WL14_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11035(__A11_NET_290, A2XG_n, A15_n, __A11_NET_291, WYHIG_n, WL15_n, GND, WL14_n, WYDG_n, __A11_NET_286, __A11_2__Y1_n, CUG, __A11_2__Y1, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11036(BXVX, __A11_NET_290, __A11_2__X1_n, CLXC, CUG, __A11_2__X1, GND, __A11_2__Y1_n, __A11_NET_291, __A11_NET_286, __A11_2__Y1, __A11_2__X1_n, __A11_2__X1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11037(__A11_NET_295, __A11_2__X1_n, __A11_2__Y1_n, __XUY15_n, __A11_2__X1, __A11_2__Y1, GND, __A11_NET_295, __XUY15_n, __A11_NET_292, __A11_NET_295, SUMA15_n, __A11_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U11038(__A11_NET_303, __A11_NET_302, SUMA15_n, SUMB15_n, RULOG_n, __A11_NET_274, GND, __A11_NET_278, XUY01_n, __XUY15_n, __CI15_n, __A11_NET_304, G15, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11039(__CI15_n, __A11_NET_293, G15_n, __A11_2___GEM1, RL15_n, WL15, GND, WL15_n, WL15,  ,  , __A11_NET_240, __A11_2___CI_INTERNAL, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11040(SUMB15_n, __A11_NET_292, __A11_NET_293, __A11_NET_277, WAG_n, WL15_n, GND, G16SW_n, WALSG_n, __A11_NET_279, A15_n, CAG, __A11_NET_275, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11041(__A11_NET_278, __A11_2___CO_OUT_U11041_2, __A11_NET_273, RL15_n_U11041_4, __A11_NET_282, L15_n_U11041_6, GND, Z15_n_U11041_8, __A11_NET_306, RL15_n_U11041_10, __A11_NET_307, RL15_n_U11041_12, __A11_NET_308, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11042(__A11_NET_277, __A11_NET_279, __A11_NET_274, __A11_NET_272, CH16, __A11_NET_273, GND, __A11_NET_282, __A11_NET_276, __A11_NET_284, __A11_NET_285, A15_n, __A11_NET_275, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11043(__A11_NET_272, RAG_n, A15_n, __A11_NET_276, WLG_n, WL15_n, GND, G01_n, G2LSG_n, __A11_NET_284, L15_n, CLG1G, __A11_NET_285, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11044(__A11_NET_242, SUMA16_n, SUMA16_n, SUMB16_n, RUG_n, __A11_NET_241, GND, __A11_2___RL_OUT_1, RLG_n, L15_n, p4VSW, EAC_n, __CO16, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11045( ,  ,  , __A11_NET_281, WQG_n, WL15_n, GND, __A11_NET_281, __A11_NET_280, __A11_2___Q1_n, __A11_2___Q1_n, CQG, __A11_NET_280, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11046(__A11_NET_283, RQG_n, __A11_2___Q1_n, __A11_NET_309, WZG_n, WL15_n, GND, __A11_NET_309, __A11_NET_310, __A11_NET_306, Z15_n, CZG, __A11_NET_310, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U11047(__A11_NET_305, RZG_n, Z15_n, __A11_NET_315, WBG_n, WL15_n, GND, __A11_NET_315, __A11_NET_314, __A11_2___B1_n, __A11_2___B1_n, CBG, __A11_NET_314, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11048(__A11_NET_312, RBHG_n, __A11_2___B1_n, __A11_NET_311, __A11_NET_314, RCG_n, GND, GND, p4VSW, __A11_NET_300, GND, p4VSW, __A11_NET_299, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11049(__A11_2___RL_OUT_1, __A11_NET_283, MDT15, R1C, __RL16, __A11_NET_308, GND, __A11_NET_313, __A11_NET_312, __A11_NET_311, __A11_NET_296, __A11_NET_307, __A11_NET_305, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11050(__A11_NET_258, __A11_2___CO_OUT_U11050_2, __A11_NET_313, RL15_n_U11050_4, __A11_NET_301, G15_n_U11050_6, GND, G15_n_U11050_8, __A11_NET_304, RL16_n_U11050_10, __A11_NET_228, L16_n_U11050_12, __A11_NET_229, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11051(__A11_NET_303, L2GDG_n, __L14_n, __A11_NET_302, WG1G_n, WL15_n, GND, G15_n, CGG, G15, RGG_n, G15_n, __A11_NET_296, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U11052(__A11_NET_301, GND, SA16, __A11_NET_300, __A11_NET_299,  , GND,  , GND, SA16, __A11_NET_264, __A11_NET_251, __A11_NET_250, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11053(__A11_NET_243, A2XG_n, A16_n, __A11_NET_247, WYHIG_n, WL16_n, GND, WL16_n, WYDG_n, __A11_NET_246, __A11_2__Y2_n, CUG, __A11_2__Y2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11054(MONEX, __A11_NET_243, __A11_2__X2_n, CLXC, CUG, __A11_2__X2, GND, __A11_2__Y2_n, __A11_NET_247, __A11_NET_246, __A11_2__Y2, __A11_2__X2_n, __A11_2__X2, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11055(__A11_NET_242, __A11_2__X2_n, __A11_2__Y2_n, __XUY16_n, __A11_2__X2, __A11_2__Y2, GND,  ,  ,  , __A11_NET_242, __XUY16_n, __A11_NET_236, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11056(SUMB16_n, __A11_NET_236, __A11_NET_240, __A11_NET_244, WAG_n, WL16_n, GND, G16SW_n, WALSG_n, __A11_NET_245, A16_n, CAG, __A11_NET_227, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U11057(__A11_NET_244, __A11_NET_245, __A11_NET_241, __A11_NET_226, CH16, __A11_NET_228, GND, __A11_NET_229, __A11_NET_263, __A11_NET_259, __A11_NET_262, A16_n, __A11_NET_227, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11058(__A11_NET_226, RAG_n, A16_n, __A11_NET_263, WLG_n, WL16_n, GND, __G16_n, G2LSG_n, __A11_NET_259, L16_n, CLG1G, __A11_NET_262, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U11059(RLG_n, L16_n, __RL16, __A11_NET_230, __A11_NET_233, __A11_NET_223, GND, __A11_NET_225, MDT16, R1C, US2SG, __RL16, GND, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11060(__A11_NET_261, WQG_n, WL16_n, __A11_2___Q2_n, __A11_NET_261, __A11_NET_231, GND, __A11_2___Q2_n, CQG, __A11_NET_231, RQG_n, __A11_2___Q2_n, __A11_NET_230, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U11061(__A11_NET_223, RL16_n_U11061_2, __A11_NET_224, Z16_n_U11061_4, __A11_NET_225, RL16_n_U11061_6, GND, RL16_n_U11061_8, __A11_NET_271, __G16_n_U11061_10, __A11_NET_250, __G16_n_U11061_12, __A11_NET_266, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11062(__A11_NET_232, WZG_n, WL16_n, __A11_NET_224, __A11_NET_232, __A11_NET_234, GND, Z16_n, CZG, __A11_NET_234, RZG_n, Z16_n, __A11_NET_233, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U11063(__A11_NET_260, WBG_n, WL16_n, __A11_2___B2_n, __A11_NET_260, __A11_NET_268, GND, __A11_2___B2_n, CBG, __A11_NET_268, RBHG_n, __A11_2___B2_n, __A11_NET_270, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U11064(__A11_NET_269, __A11_NET_268, RCG_n, __A11_NET_264, WL14_n, WG3G_n, GND, WL01_n, WG5G_n, __A11_NET_251, L2GDG_n, L16_n, __A11_NET_265, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U11065(__G16_n, GEM16, RL16_n, WL16, WL16, WL16_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U11066(SUMA13_n, __A11_NET_202, XUY13_n, CI13_n, GND,  , GND,  , __A11_NET_148, XUY14_n, __A11_1___CI_INTERNAL, GND, SUMA14_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U11067(SUMA15_n, __A11_NET_295, __XUY15_n, __CI15_n, GND,  , GND,  , __A11_NET_242, __XUY16_n, __A11_2___CI_INTERNAL, WHOMPA, SUMA16_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U11068(RL13_n, MWL13_U11068_2, RL14_n, MWL14_U11068_4, RL15_n, MWL15_U11068_6, GND, MWL16_U11068_8, RL16_n,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12001(G01, __A12_1__G01A_n, G02, __A12_1__G02_n, G03, __A12_1__G03_n, GND, __A12_1__PA03_n, __A12_1__PA03, __A12_NET_184, G04, __A12_NET_183, G05, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12002(G01, G02, G01, __A12_1__G02_n, __A12_1__G03_n, __A12_NET_178, GND, __A12_NET_179, __A12_1__G01A_n, G02, __A12_1__G03_n, __A12_NET_206, G03, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12003(__A12_1__G01A_n, __A12_1__G02_n, G04, G05, G06, __A12_NET_200, GND, __A12_NET_198, G04, __A12_NET_183, __A12_NET_187, __A12_NET_180, G03, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U12004(__A12_1__PA03, __A12_NET_206, __A12_NET_178, __A12_NET_179, __A12_NET_180,  , GND,  , __A12_NET_200, __A12_NET_198, __A12_NET_185, __A12_NET_195, __A12_1__PA06, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12005(G06, __A12_NET_187, __A12_NET_200, __A12_NET_136, __A12_1__PA06, __A12_1__PA06_n, GND, __A12_NET_188, G07, __A12_NET_199, G08, __A12_NET_189, G09, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12006(__A12_NET_184, G05, __A12_NET_184, __A12_NET_183, G06, __A12_NET_195, GND, __A12_NET_201, G07, G08, G09, __A12_NET_185, __A12_NET_187, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12007(G07, __A12_NET_199, __A12_NET_188, G08, __A12_NET_189, __A12_NET_190, GND, __A12_NET_191, __A12_NET_188, __A12_NET_199, G09, __A12_NET_192, __A12_NET_189, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U12008(__A12_1__PA09, __A12_NET_201, __A12_NET_192, __A12_NET_190, __A12_NET_191,  , GND,  , __A12_NET_126, __A12_NET_123, __A12_NET_124, __A12_NET_125, __A12_1__PA12, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12009(__A12_NET_201, __A12_NET_137, __A12_1__PA09, __A12_1__PA09_n, G10, __A12_NET_168, GND, __A12_NET_122, G11, __A12_NET_167, G12, __A12_NET_128, __A12_NET_126, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12010(G10, G11, G10, __A12_NET_122, __A12_NET_167, __A12_NET_123, GND, __A12_NET_124, __A12_NET_168, G11, __A12_NET_167, __A12_NET_126, G12, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12011(__A12_NET_168, __A12_NET_122, G13, G14, G16, __A12_NET_135, GND, __A12_NET_132, G13, __A12_NET_121, __A12_1__G16A_n, __A12_NET_125, G12, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12012(__A12_1__PA12, __A12_1__PA12_n, G13, __A12_NET_127, G14, __A12_NET_121, GND, __A12_1__G16A_n, G16, __A12_NET_129, __A12_NET_135, __A12_1__PA15_n, __A12_1__PA15, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12013(__A12_NET_127, G14, __A12_NET_127, __A12_NET_121, G16, __A12_NET_134, GND, __A12_NET_173, __A12_NET_136, __A12_NET_137, __A12_NET_128, __A12_NET_133, __A12_1__G16A_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U12014(__A12_1__PA15, __A12_NET_135, __A12_NET_132, __A12_NET_133, __A12_NET_134,  , GND,  , EXTPLS, RELPLS, INHPLS, __A12_NET_119, __A12_NET_118, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12015(__A12_NET_171, __A12_NET_129, G15, __A12_NET_131, TSUDO_n, __A12_1__T7PHS4_n, GND, __A12_1__G02_n, G03, __A12_NET_204, G02, __A12_1__G03_n, __A12_NET_203, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U12016(__A12_NET_173, __A12_1__GNZRO_U12016_2, __A12_NET_171, __A12_1__GNZRO_U12016_4, __A12_NET_205, RELPLS_U12016_6, GND, RELPLS_U12016_8, __A12_NET_204, INHPLS_U12016_10, __A12_NET_202, INHPLS_U12016_12, __A12_NET_203, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12017(__A12_1__GNZRO, __A12_NET_113, __A12_NET_178, __A12_NET_130, __A12_NET_131, __A12_NET_114, GND, GEQZRO_n, __A12_NET_112, __A12_NET_120, RAD, __A12_1__PB09_n, __A12_1__PB09, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12018(__A12_NET_130, __A12_NET_113, __A12_NET_113, __A12_NET_114, __A12_1__G01A_n, __A12_NET_205, GND, __A12_NET_202, __A12_NET_113, G01, __A12_NET_114, EXTPLS, __A12_NET_114, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U12019(__A12_NET_112, __A12_NET_113, G02, G01, G03,  , GND,  , __A12_NET_162, __A12_NET_115, __A12_NET_117, __A12_NET_153, __A12_1__PB09, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12020(__A12_NET_119, __A12_NET_118, T12A, RADRZ, __A12_NET_118, __A12_NET_120, GND, __A12_NET_120, __A12_NET_119, RADRG, __A12_1__PA12, __A12_1__PA15, __A12_NET_151, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12021(__A12_1__PA03, __A12_1__PA06, __A12_1__PA03, __A12_1__PA06_n, __A12_1__PA09_n, __A12_NET_115, GND, __A12_NET_117, __A12_1__PA03_n, __A12_1__PA06, __A12_1__PA09_n, __A12_NET_162, __A12_1__PA09, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U12022(__A12_1__PA03_n, __A12_1__PA06_n, __A12_NET_142, MONPAR, SAP, __A12_NET_143, GND, __A12_NET_139, SCAD, __A12_NET_140, GOJAM, __A12_NET_153, __A12_1__PA09, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12023(__A12_NET_149, __A12_1__PA12_n, __A12_1__PA15_n, __A12_1__PB15, __A12_NET_151, __A12_NET_149, GND, __A12_1__PB09_n, __A12_1__PB15, __A12_NET_160, __A12_1__PB09, __A12_1__PB15_n, __A12_NET_161, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12024(__A12_1__PB15, __A12_1__PB15_n, __A12_1__PC15, PC15_n, __A12_1__PC15, MGP_n, GND, GEMP, PC15_n, MSP, __A12_NET_143,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12025(__A12_1__PC15, __A12_NET_160, __A12_NET_161, __A12_NET_142, CGG, __A12_NET_143, GND, __A12_1__PC15, __A12_NET_142, __A12_NET_140, PC15_n, __A12_NET_143, __A12_NET_138, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12026(TPARG_n, n8XP5, T07_n, PHS4_n, FUTEXT, __A12_1__T7PHS4, GND, __A12_NET_231, XB0_n, T02_n, __A12_NET_233, __A12_NET_141, __A12_NET_138, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U12027(__A12_NET_139, PALE_U12027_2, __A12_NET_141, PALE_U12027_4,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12028(G01ED, WEDOPG_n, WL08_n, __A12_NET_249, WL08_n, WSG_n, GND, __A12_NET_249, __A12_NET_250, __A12_NET_251, __A12_NET_251, CSG, __A12_NET_250, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12029(__A12_NET_251, S08, __A12_NET_250, S08_n, __A12_NET_247, S09, GND, S09_n, __A12_NET_248, S10, __A12_NET_256, S10_n, __A12_NET_257, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12030(G02ED, WEDOPG_n, WL09_n, __A12_NET_246, WL09_n, WSG_n, GND, __A12_NET_246, __A12_NET_248, __A12_NET_247, __A12_NET_247, CSG, __A12_NET_248, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12031(G03ED, WEDOPG_n, WL10_n, __A12_NET_255, WL10_n, WSG_n, GND, __A12_NET_255, __A12_NET_257, __A12_NET_256, __A12_NET_256, CSG, __A12_NET_257, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12032(G04ED, WEDOPG_n, WL11_n, __A12_NET_252, WL11_n, WSG_n, GND, __A12_NET_252, __A12_NET_254, __A12_NET_253, __A12_NET_253, CSG, __A12_NET_254, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12033(__A12_NET_253, S11, __A12_NET_254, S11_n, __A12_NET_244, S12, GND, S12_n, __A12_NET_245, S01, __A12_NET_219, S01_n, __A12_NET_218, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12034(G05ED, WEDOPG_n, WL12_n, __A12_NET_243, WL12_n, WSG_n, GND, EDOP_n, T12A, __A12_NET_239, __A12_NET_244, CSG, __A12_NET_245, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U12035(G06ED, WEDOPG_n, WL13_n, G07ED, WEDOPG_n, WL14_n, GND, WL01_n, WSG_n, __A12_NET_225, __A12_NET_225, __A12_NET_218, __A12_NET_219, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12036(__A12_NET_218, __A12_NET_219, CSG, __A12_NET_226, WL02_n, WSG_n, GND, __A12_NET_226, __A12_NET_216, __A12_NET_217, __A12_NET_217, CSG, __A12_NET_216, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12037(__A12_NET_217, S02, __A12_NET_216, S02_n, __A12_NET_215, S03, GND, S03_n, __A12_NET_214, S04, __A12_NET_213, S04_n, __A12_NET_227, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U12038(__A12_NET_229, WL03_n, WSG_n, __A12_NET_215, __A12_NET_229, __A12_NET_214, GND, __A12_NET_215, CSG, __A12_NET_214, WL04_n, WSG_n, __A12_NET_230, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U12039(__A12_NET_213, __A12_NET_230, __A12_NET_227, __A12_NET_227, __A12_NET_213, CSG, GND, WL05_n, WSG_n, __A12_NET_228, __A12_NET_228, __A12_NET_211, __A12_NET_212, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U12040(__A12_NET_211, __A12_NET_212, CSG, __A12_NET_220, WL06_n, WSG_n, GND, __A12_NET_220, __A12_NET_209, __A12_NET_210, __A12_NET_210, CSG, __A12_NET_209, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12041(__A12_NET_212, S05, __A12_NET_211, S05_n, __A12_NET_210, S06, GND, S06_n, __A12_NET_209, S07, __A12_NET_208, S07_n, __A12_NET_207, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U12042(__A12_NET_221, WL07_n, WSG_n, __A12_NET_208, __A12_NET_221, __A12_NET_207, GND, __A12_NET_208, CSG, __A12_NET_207,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U12043(__A12_1__T7PHS4, __A12_1__T7PHS4_n,  ,  , OCTAD2, __A12_NET_233, GND, GINH, __A12_NET_222, __A12_2__G01A, __A12_1__G01A_n,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U12044( ,  ,  ,  ,  ,  , GND,  , __A12_NET_223, __A12_NET_232, __A12_NET_240, __A12_NET_239, __A12_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U12045( ,  ,  , CYR_n, __A12_NET_231, __A12_NET_223, GND, CYR_n, T12A, __A12_NET_223, __A12_NET_234, __A12_NET_232, SR_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U12046(__A12_NET_233, T02_n, __A12_NET_233, T02_n, XB2_n, __A12_NET_241, GND, __A12_NET_238, __A12_NET_233, T02_n, XB3_n, __A12_NET_234, XB1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U12047(__A12_NET_232, SR_n, T12A, CYL_n, __A12_NET_241, __A12_NET_240, GND, CYL_n, T12A, __A12_NET_240, __A12_NET_238, __A12_NET_239, EDOP_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U12048(n8XP5, __A12_NET_243, SUMA16_n, SUMB16_n, __A12_1__G01A_n, __A12_NET_237, GND,  ,  ,  ,  , __A12_NET_244, __A12_NET_245, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U12049(__A12_NET_236, __A12_2__G01A, __A12_1__G16A_n, G16SW_n, __A12_NET_236, __A12_NET_237, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U12050(PALE, MPAL_n_U12050_2,  ,  ,  ,  ,  ,  ,  ,  ,  ,  ,  ,  , SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U13001(MSTRT, __A13_NET_255, F12B, __A13_1__F12B_n, __A13_1__F14H, __A13_NET_242, GND, __A13_NET_274, __A13_NET_277, __A13_1__NOTEST, __A13_1__NOTEST_n, __A13_1__DOFILT, __A13_NET_264, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13002(__A13_NET_254, F05B_n, __A13_NET_255, __A13_NET_253, __A13_NET_254, __A13_NET_201, GND, __A13_NET_253, __A13_NET_255, __A13_NET_201, F05A_n, __A13_NET_253, MSTRTP, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U13003(__A13_NET_257, IIP, __A13_NET_256, __A13_NET_256, __A13_NET_257, F14B, GND, IIP_n, __A13_NET_241, __A13_NET_238, __A13_NET_238, F14B, __A13_NET_241, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13004(__A13_1__F12B_n, FS14, PALE, __A13_NET_243, __A13_NET_235, __A13_NET_251, GND, __A13_NET_252, __A13_NET_248, __A13_NET_237, __A13_1__WATCHP, __A13_1__F14H, __A13_1__FS13_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U13005(__A13_NET_243, __A13_NET_256, __A13_NET_242, __A13_NET_235, __A13_NET_241, __A13_NET_242, GND, __A13_NET_243, __A13_NET_235, __A13_NET_205, __A13_NET_234, F10B, __A13_NET_233, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U13006(__A13_NET_251, __A13_1__CKTAL_n_U13006_2, __A13_NET_252, __A13_1__CKTAL_n_U13006_4, __A13_NET_227, __A13_NET_277_U13006_6, GND, __A13_NET_277_U13006_8, __A13_NET_228, __A13_NET_277_U13006_10, __A13_NET_220, __A13_NET_277_U13006_12, __A13_NET_221, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U13007(TC0, TCF0, T12_n, PHS4_n, NISQL_n, __A13_NET_309, GND, __A13_NET_281, __A13_1__NOTEST, __A13_NET_272, T09_n, __A13_NET_234, __A13_NET_233, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13008(__A13_NET_231, __A13_NET_236, __A13_NET_232, __A13_NET_232, __A13_NET_231, F10B, GND, __A13_NET_233, F10A_n, __A13_NET_248, __A13_NET_232, F10A_n, __A13_NET_237, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U13009(__A13_NET_236, TCF0, TC0, INKL, T04_n,  , GND,  , INLNKP, INLNKM, RNRADP, RNRADM, __A13_NET_196, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13010(__A13_NET_206, __A13_NET_248, __A13_NET_237, __A13_NET_272, __A13_NET_274, __A13_NET_273, GND, __A13_NET_272, INKL, __A13_NET_273, PSEUDO, NISQL_n, __A13_1__NOTEST_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U13011(__A13_NET_197, GYROD, CDUXD, CDUYD, CDUZD,  , GND,  , TRUND, SHAFTD, THRSTD, EMSD, __A13_NET_198, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13012(__A13_NET_284, __A13_NET_281, __A13_NET_282, __A13_NET_282, __A13_NET_284, INKL, GND, T03_n, __A13_NET_284, __A13_NET_283, __A13_NET_283, __A13_NET_262, __A13_NET_207, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13013(INKL, T03_n, __A13_NET_283, __A13_NET_262, GOJAM, __A13_NET_264, GND, __A13_NET_315, __A13_NET_313, __A13_NET_314, __A13_NET_304, __A13_NET_279, CTROR, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13014(__A13_NET_278, __A13_NET_279, __A13_NET_280, __A13_NET_280, __A13_NET_278, F07A, GND, __A13_NET_280, F07B_n, __A13_NET_262, NHALGA, __A13_1__CKTAL_n, ALGA, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U13115(__A13_1__SCAS10, __A13_1__CON2, FS10, __A13_1__SCAS17, FS17, DOSCAL, GND, F05B_n, __A13_NET_266, __A13_NET_261, __A13_NET_261, __A13_NET_260, __A13_NET_267, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U13116(VFAIL, __A13_NET_266,  ,  , TEMPIN, __A13_1__TEMPIN_n, GND,  ,  , __A13_NET_178, F14B, __A13_1__FILTIN, __A13_NET_189, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U13117(__A13_NET_267, __A13_NET_266, F05A_n, __A13_NET_267, NHVFAL, __A13_NET_204, GND, __A13_NET_268, F05A_n, __A13_NET_267, STNDBY_n, __A13_NET_260, NHVFAL, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13118(__A13_NET_270, __A13_NET_204, STRT1, STRT1, __A13_NET_270, __A13_NET_271, GND, __A13_NET_260, F05A_n, __A13_NET_271, __A13_1__CON3, n2FSFAL, __A13_1__SCADBL, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U13119(__A13_NET_268, __A13_1__DOFILT, SB0_n, __A13_NET_179, __A13_NET_178, __A13_NET_180, GND, __A13_NET_187, FLTOUT, SCAFAL, AGCWAR, __A13_NET_183, __A13_1__SCADBL, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U13120(__A13_1__CON3, __A13_1__CON2, FS10,  ,  ,  , GND, ALTEST, __A13_NET_184, __A13_NET_177, __A13_NET_179, __A13_NET_176, __A13_NET_184, p4VDC, SIM_RST, SIM_CLK);
    U74LVC07 U13121(__A13_NET_183, __A13_NET_179_U13121_2, __A13_NET_177, __A13_NET_179_U13121_4,  ,  , GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13122(__A13_NET_176, SB2_n, __A13_NET_178, __A13_NET_189, __A13_NET_180, __A13_NET_188, GND, __A13_NET_189, F08B, __A13_NET_188, FLTOUT, SCAFAL, __A13_NET_186, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U13123(__A13_NET_186, __A13_1__WARN, __A13_1__WARN, __A13_1__CGCWAR,  ,  , GND,  ,  ,  ,  , TMPCAU, __A13_NET_164, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U13124(AGCWAR, __A13_NET_187, CCH33, __A13_NET_167, STRT2, OSCALM, GND, __A13_NET_167, CCH33, OSCALM, __A13_1__TEMPIN_n, TMPOUT, __A13_NET_164, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U13125(__A13_NET_166, GOJAM, __A13_NET_165, __A13_NET_172, ALTEST, __A13_NET_165, GND, SBY, __A13_NET_174, __A13_NET_175, __A13_NET_175, T10, __A13_NET_174, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U13126(__A13_NET_166, ERRST, CT_n, P02_n, P03, __A13_NET_170, GND,  ,  ,  ,  , __A13_NET_165, __A13_1__SBYEXT, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U13127(__A13_NET_172, RESTRT, __A13_NET_175, __A13_1__SBYEXT, __A13_NET_171, __A13_1__SYNC4_n, GND, __A13_1__SYNC14_n, __A13_NET_170,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC4002 U13128(__A13_NET_171, FS01, P02, P03_n, CT_n,  , GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U13029(__A13_NET_217, __A13_NET_215, __A13_NET_216, __A13_NET_216, __A13_NET_217, F17B, GND, __A13_NET_211, SB1_n, __A13_NET_212, __A13_1__WATCHP, __A13_1__WATCH, __A13_NET_213, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13030(SB2_n, __A13_NET_216, __A13_NET_313, __A13_NET_310, __A13_NET_304, __A13_NET_321, GND, __A13_NET_312, __A13_NET_313, __A13_NET_311, __A13_NET_304, __A13_1__WATCHP, __A13_NET_211, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b1) U13031(__A13_1__WATCH, __A13_NET_213, __A13_NET_212, __A13_NET_190, OTLNKM, ALTM, GND, __A13_NET_306, __A13_NET_305, __A13_NET_304, __A13_NET_315, __A13_NET_323, __A13_NET_322, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U13032( ,  , __A13_NET_307, __A13_NET_313, MLOAD, __A13_NET_314, GND, __A13_NET_310, MREAD, __A13_NET_311, MLDCH, __A13_NET_302, MRDCH, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U13033(__A13_NET_228, T5P, T6P, CDUXP, CDUXM,  , GND,  , CDUYP, CDUYM, CDUZP, CDUZM, __A13_NET_220, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U13034(__A13_NET_221, TRNP, TRNM, SHAFTP, SHAFTM,  , GND,  , PIPXP, PIPXM, PIPYP, PIPYM, __A13_NET_191, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U13035(__A13_NET_195, PIPZP, PIPZM, BMAGXP, BMAGXM,  , GND,  , BMAGYP, BMAGYM, BMAGZP, BMAGZM, __A13_NET_192, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U13036(__A13_NET_197, __A13_NET_277_U13036_2, __A13_NET_198, __A13_NET_277_U13036_4, __A13_NET_190, __A13_NET_277_U13036_6, GND, __A13_NET_307_U13036_8, __A13_NET_309, __A13_NET_307_U13036_10, __A13_NET_308, __A13_NET_277_U13036_12, __A13_NET_191, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13037(__A13_NET_313, __A13_NET_302, __A13_NET_304, GOJAM, __A13_NET_287, __A13_NET_305, GND, __A13_NET_323, __A13_NET_322, GOJAM, __A13_NET_318, __A13_NET_303, __A13_NET_304, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U13038(__A13_NET_301, MRDCH, MLDCH, MREAD, MLOAD,  , GND,  , __A13_NET_323, __A13_NET_320, INOTLD, __A13_2__INOTRD, __A13_NET_286, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b1) U13039(__A13_NET_319, __A13_NET_321, __A13_NET_320, __A13_NET_324, __A13_NET_312, INOTLD, GND, __A13_NET_324, __A13_NET_316, INOTLD, __A13_NET_303, __A13_2__INOTRD, __A13_NET_317, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13040(__A13_NET_319, GOJAM, MON_n, __A13_NET_290, ST1_n, __A13_NET_318, GND, __A13_NET_316, T12_n, CT, PHS2_n, __A13_NET_320, __A13_NET_318, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U13041(__A13_2__INOTRD, __A13_NET_317, __A13_NET_316, __A13_2__STORE1, ST1_n, __A13_NET_322, GND, ST1_n, __A13_NET_319, FETCH1, __A13_NET_323, __A13_NET_320, MON_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U13042(FETCH0, ST0_n, MON_n, STFET1_n, __A13_2__STORE1, FETCH1, GND, __A13_NET_285, T11_n, __A13_NET_287, CTROR_n, __A13_NET_305, __A13_NET_294, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U13043(__A13_NET_316, __A13_NET_290, __A13_2__STORE1, STORE1_n, FETCH0, FETCH0_n, GND, MONpCH, __A13_NET_286,  ,  , INCSET_n, __A13_NET_297, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13044(FETCH1, __A13_2__STORE1, __A13_NET_294, T12_n, PHS3_n, __A13_NET_295, GND, __A13_NET_292, __A13_NET_291, __A13_NET_295, GOJAM, __A13_NET_285, CHINC, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U13045(__A13_NET_293, __A13_NET_313, MNHNC, __A13_NET_305, CTROR_n,  , GND,  , T1P, T2P, T3P, T4P, __A13_NET_227, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U13046(__A13_NET_291, __A13_NET_293, __A13_NET_292, __A13_NET_297, T02_n, __A13_NET_291, GND, __A13_NET_292, MONpCH, INKL_n, __A13_2__INOTRD, INOTLD, CHINC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U13047(INKL_n, INKL,  ,  , T10_n, BKTF_n, GND, CHINC, CHINC_n, __A13_1__FS13_n, FS13, __A13_1__CON1, DBLTST, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U13048(__A13_NET_291, T07_n, T02_n, CA6_n, XB7_n, __A13_NET_215, GND,  ,  ,  ,  , RSSB, PHS3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U13049(__A13_NET_308, GNHNC, PSEUDO, __A13_NET_306, PHS2_n, __A13_NET_301, GND, __A13_1__CON1, FS09, __A13_1__CON2,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U13050( ,  ,  ,  ,  ,  , GND,  ,  ,  ,  , __A13_NET_211, F17A, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U13051(__A13_NET_195, __A13_NET_277_U13051_2, __A13_NET_192, __A13_NET_277_U13051_4, __A13_NET_196, __A13_NET_277_U13051_6, GND, MRPTAL_n_U13051_8, __A13_NET_205, MTCAL_n_U13051_10, __A13_NET_206, MCTRAL_n_U13051_12, __A13_NET_207, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U13052(__A13_NET_204, MVFAIL_n_U13052_2, PIPAFL, MPIPAL_n_U13052_4, __A13_1__SCADBL, MSCDBL_n_U13052_6, GND, MWATCH_n_U13052_8, __A13_1__WATCH, MSCAFL_n_U13052_10, SCAFAL, MWARNF_n_U13052_12, FLTOUT, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U13053(STRT2, MOSCAL_n_U13053_2, INKL_n, MINKL_U13053_4, __A13_NET_286, MREQIN_U13053_6, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U14001(__A14_1__ROP_n, S11, S12, __A14_NET_192, T08_n, PHS3_n, GND, __A14_NET_192, __A14_NET_193, __A14_NET_202, __A14_NET_201, __A14_NET_198, __A14_NET_200, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14002(__A14_NET_202, T09, __A14_1__ROP_n, __A14_NET_202, T08, __A14_NET_201, GND, __A14_NET_198, __A14_NET_200, __A14_NET_231, TIMR, __A14_NET_193, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14003(T01_n, __A14_NET_231, __A14_NET_200, __A14_1__IHENV, __A14_NET_228, __A14_1__SETAB_n, GND, SETAB, __A14_1__SETAB_n, __A14_1__SETCD_n, __A14_NET_227, SETCD, __A14_1__SETCD_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14004(TIMR, __A14_NET_231, PHS4_n, __A14_1__ROP_n, T10_n, __A14_NET_230, GND, __A14_NET_237, T05_n, PHS3_n, __A14_1__ROP_n, __A14_NET_199, __A14_NET_229, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14005(__A14_NET_229, __A14_NET_199, __A14_NET_230, __A14_NET_228, S09, __A14_NET_229, GND, __A14_NET_229, S09_n, __A14_NET_227, __A14_NET_237, __A14_NET_236, __A14_NET_235, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14006(__A14_NET_235, T08, __A14_NET_235, S09, S08, __A14_NET_234, GND, __A14_NET_232, __A14_NET_235, S09, S08_n, __A14_NET_236, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U14007(__A14_NET_233, __A14_1__CLEARA, __A14_NET_234, __A14_NET_224, __A14_1__CLEARB, __A14_NET_232, GND, __A14_1__CLEARC, __A14_NET_221, __A14_NET_220, __A14_1__CLEARD, __A14_NET_217, __A14_NET_219, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14008(__A14_NET_233, RESETA, __A14_NET_224, RESETB, __A14_NET_220, RESETC, GND, RESETD, __A14_NET_219, __A14_1__S08A_n, S08, __A14_1__S08A, S08_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14009(__A14_NET_235, S08, __A14_NET_235, S09_n, S08_n, __A14_NET_217, GND, STBF, GOJAM, __A14_NET_223, __A14_NET_269, __A14_NET_221, S09_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U14010(__A14_1__CLEARA, __A14_1__SETAB_n, __A14_1__S08A_n, __A14_1__CLEARB, __A14_1__SETAB_n, __A14_1__S08A, GND, __A14_1__SETCD_n, __A14_1__S08A_n, __A14_1__CLEARC, __A14_1__SETCD_n, __A14_1__S08A, __A14_1__CLEARD, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14011(__A14_NET_269, STBF, __A14_1__SBFSET, __A14_NET_223, T07_n, PHS3_n, GND, T02_n, __A14_1__ROP_n, __A14_NET_280, __A14_NET_280, STRGAT, __A14_NET_274, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14012(__A14_NET_269, SBF, __A14_1__ROP_n, __A14_NET_194, S07_n, __A14_2__IL07_n, GND, WEX, __A14_NET_206, WEY, __A14_NET_203, __A14_1__ERAS_n, __A14_1__ERAS, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14013(MNHSBF, MP1, __A14_1__ROP_n, T06_n, DV3764, __A14_NET_270, GND, STRGAT, __A14_NET_274, T08, GOJAM, __A14_NET_268, PHS4_n, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U14014(__A14_NET_268, __A14_1__SBFSET_U14014_2, __A14_NET_270, __A14_1__SBFSET_U14014_4, __A14_NET_273, __A14_1__TPGF_U14014_6, GND, __A14_1__TPGF_U14014_8, __A14_NET_279, __A14_1__ERAS_U14014_10, __A14_NET_286, __A14_1__ERAS_U14014_12, __A14_NET_285, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U14015(__A14_NET_273, __A14_1__ROP_n, T08_n, DV3764, GOJ1,  , GND,  , GOJAM, TCSAJ3, PHS2_n, MP1, __A14_NET_279, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14016(T02_n, __A14_NET_194, __A14_NET_196, T03, GOJAM, __A14_NET_197, GND, __A14_NET_213, __A14_NET_211, T07, GOJAM, __A14_NET_212, __A14_NET_196, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U14017(__A14_NET_195, __A14_1__ROP_n, T10_n, __A14_NET_196, __A14_NET_195, __A14_NET_197, GND, __A14_NET_212, __A14_NET_213, __A14_NET_211, T01, __A14_NET_214, __A14_NET_215, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14018(__A14_NET_214, __A14_NET_215, __A14_NET_216, __A14_NET_216, T12_n, PHS3_n, GND, T12A, __A14_NET_214, __A14_NET_207, __A14_NET_205, __A14_NET_210, __A14_NET_206, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14019(__A14_NET_207, TIMR, __A14_NET_207, TIMR, __A14_NET_203, __A14_NET_204, GND, __A14_NET_209, TIMR, T11, __A14_NET_208, __A14_NET_205, __A14_NET_206, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b0) U14020(__A14_NET_203, __A14_NET_204, __A14_NET_251, __A14_NET_208, __A14_NET_209, __A14_NET_252, GND, __A14_NET_208, T10, __A14_NET_210, T05_n, __A14_1__ERAS_n, __A14_NET_256, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14021(__A14_NET_259, __A14_NET_260, __A14_1__ERAS_n, PHS3_n, T03_n, __A14_NET_261, GND, __A14_NET_257, __A14_1__FNERAS_n, T12A, GOJAM, __A14_NET_258, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U14022(__A14_1__FNERAS_n, __A14_NET_256, __A14_NET_257, __A14_NET_266, __A14_1__FNERAS_n, T10_n, GND, __A14_NET_254, __A14_NET_252, __A14_NET_253, T02_n, PHS4_n, __A14_NET_263, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14023(T10_n, __A14_1__FNERAS_n, __A14_1__FNERAS_n, T10_n, PHS3_n, __A14_NET_252, GND, __A14_NET_254, TIMR, __A14_NET_263, __A14_NET_253, __A14_NET_251, PHS4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14024(TIMR, T01, __A14_NET_241, GOJAM, __A14_1__REDRST, __A14_NET_262, GND, __A14_NET_243, __A14_NET_242, GOJAM, __A14_1__REDRST, __A14_NET_265, __A14_NET_264, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U14025(__A14_NET_264, __A14_NET_265, __A14_NET_266, ZID, __A14_NET_264, MYCLMP, GND, __A14_1__ERAS_n, T03_n, __A14_NET_267, __A14_NET_267, __A14_NET_258, __A14_NET_259, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U14026(__A14_NET_286, TCSAJ3, S11, S12, INOUT,  , GND,  , CHINC, GOJ1, MP1, MAMU, __A14_NET_285, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b1) U14027(SETEK, MYCLMP, __A14_NET_259, __A14_NET_260, T06_n, PHS3_n, GND, __A14_NET_261, __A14_NET_262, __A14_NET_241, __A14_NET_244, __A14_NET_243, __A14_NET_242, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14028(__A14_NET_241, REY, __A14_NET_242, REX, __A14_NET_238, SBE, GND, __A14_1__RSTK_n, __A14_NET_253, RSTKY_n, __A14_1__RSTK_n, RSTKX_n, __A14_1__RSTK_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14029(__A14_1__ERAS_n, T03_n, GOJAM, T05, __A14_NET_238, STBE, GND, __A14_1__SBESET, T04_n, __A14_1__ERAS_n, SCAD, __A14_NET_244, PHS4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U14030(__A14_1__REDRST, __A14_NET_245, T05, __A14_NET_245, __A14_NET_239, __A14_NET_240, GND, __A14_NET_245, T06, __A14_NET_240, T05_n, PHS3_n, __A14_NET_239, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U14031(__A14_NET_238, STBE, __A14_1__SBESET, __A14_NET_249, T05_n, PHS3_n, GND, __A14_1__TPGF, __A14_1__TPGE, TPARG_n, S07, S08, __A14_2__YB0, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14032(SCAD, __A14_1__ERAS_n, S01, S02, S03, XB0, GND, XB1, S01_n, S02, S03, __A14_NET_248, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U14033(__A14_NET_248, __A14_1__TPGE_U14033_2, __A14_NET_249, __A14_1__TPGE_U14033_4,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14034(XB0, XB0_n, XB0_n, __A14_2__XB0E, XB1, XB1_n, GND, XB1E, XB1_n, XB2_n, XB2, XB2E, XB2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14035(S01, S02_n, S01_n, S02_n, S03, XB3, GND, XB4, S01, S02, S03_n, XB2, S03, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14036(XB3, XB3_n, XB3_n, XB3E, XB4, XB4_n, GND, XB4E, XB4_n, XB5_n, XB5, XB5E, XB5_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14037(S01_n, S02, S01, S02_n, S03_n, XB6, GND, XB7, S01_n, S02_n, S03_n, XB5, S03_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14038(XB6, XB6_n, XB6_n, XB6E, XB7, XB7_n, GND, XB7E, XB7_n, YB0_n, __A14_2__YB0, __A14_2__YB0E, YB0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U14039(__A14_2__YB1, S07_n, S08, __A14_2__YB2, S07, S08_n, GND, S07_n, S08_n, __A14_2__YB3, EB9, S10_n, __A14_NET_290, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14040(__A14_2__YB1, __A14_2__YB1_n, __A14_2__YB1_n, YB1E, __A14_2__YB2, __A14_2__YB2_n, GND, YB2E, __A14_2__YB2_n, __A14_2__YB3_n, __A14_2__YB3, YB3E, __A14_2__YB3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14041(S04, S05, S04_n, S05, S06, __A14_2__XT1, GND, __A14_2__XT2, S04, S05_n, S06, __A14_2__XT0, S06, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14042(__A14_2__XT0, XT0_n, XT0_n, __A14_2__XT0E, __A14_2__XT1, XT1_n, GND, XT1E, XT1_n, XT2_n, __A14_2__XT2, XT2E, XT2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14043(S04_n, S05_n, S04, S05, S06_n, __A14_2__XT4, GND, __A14_2__XT5, S04_n, S05, S06_n, __A14_2__XT3, S06, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14044(__A14_2__XT3, XT3_n, XT3_n, XT3E, __A14_2__XT4, XT4_n, GND, XT4E, XT4_n, XT5_n, __A14_2__XT5, XT5E, XT5_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14045(S04, S05_n, S04_n, S05_n, S06_n, __A14_2__XT7, GND, __A14_2__EAD11, S09_n, S10_n, EB11_n, __A14_2__XT6, S06_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14046(__A14_2__XT6, XT6_n, XT6_n, XT6E, __A14_2__XT7, __A14_2__XT7_n, GND, XT7E, __A14_2__XT7_n, __A14_2__EAD09_n, __A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD10, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U14047(__A14_2__EAD09, __A14_NET_290, S09_n, __A14_NET_291, EB10, S09_n, GND, S10_n, __A14_NET_291, __A14_2__EAD10, __A14_2__YB0, __A14_2__YB3, __A14_2__RILP1, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14048(__A14_2__EAD11, __A14_2__EAD11_n, __A14_2__YT0, YT0_n, YT0_n, __A14_2__YT0E, GND, __A14_2__YT1_n, __A14_2__YT1, YT1E, __A14_2__YT1_n, __A14_2__YT2_n, __A14_2__YT2, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14049(__A14_2__EAD09, __A14_2__EAD10, __A14_2__EAD09_n, __A14_2__EAD10, __A14_2__EAD11, __A14_2__YT1, GND, __A14_2__YT2, __A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD11, __A14_2__YT0, __A14_2__EAD11, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14050(__A14_2__YT2_n, YT2E, __A14_2__YT3, __A14_2__YT3_n, __A14_2__YT3_n, YT3E, GND, __A14_2__YT4_n, __A14_2__YT4, YT4E, __A14_2__YT4_n, __A14_2__YT5_n, __A14_2__YT5, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14051(__A14_2__EAD09_n, __A14_2__EAD10_n, __A14_2__EAD09, __A14_2__EAD10, __A14_2__EAD11_n, __A14_2__YT4, GND, __A14_2__YT5, __A14_2__EAD09_n, __A14_2__EAD10, __A14_2__EAD11_n, __A14_2__YT3, __A14_2__EAD11, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14052(__A14_2__YT5_n, YT5E, __A14_2__YT6, __A14_2__YT6_n, __A14_2__YT6_n, YT6E, GND, __A14_2__YT7_n, __A14_2__YT7, YT7E, __A14_2__YT7_n, __A14_NET_305, __A14_NET_302, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14053(__A14_2__EAD09, __A14_2__EAD10_n, __A14_2__EAD09_n, __A14_2__EAD10_n, __A14_2__EAD11_n, __A14_2__YT7, GND, __A14_NET_296, __A14_NET_302, __A14_2__RILP1, __A14_NET_301, __A14_2__YT6, __A14_2__EAD11_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U14054(__A14_NET_302, XB0, XB3, XB5, XB6,  , GND,  , __A14_2__XT0, __A14_2__XT3, __A14_2__XT5, __A14_2__XT6, __A14_NET_301, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14055(__A14_NET_301, __A14_NET_294, __A14_2__RILP1, __A14_2__RILP1_n, __A14_NET_295, __A14_NET_292, GND, __A14_2__ILP_n, __A14_NET_295, __A14_2__ILP, __A14_NET_292, IL01, S01, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U14056(__A14_NET_305, __A14_2__RILP1, __A14_NET_305, __A14_2__RILP1_n, __A14_NET_301, __A14_NET_299, GND, __A14_NET_300, __A14_NET_302, __A14_2__RILP1_n, __A14_NET_294, __A14_NET_298, __A14_NET_294, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U14057(__A14_NET_295, __A14_NET_296, __A14_NET_298, __A14_NET_299, __A14_NET_300,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14058(S01_n, __A14_2__IL01_n, S02, IL02, S02_n, __A14_2__IL02_n, GND, IL03, S03, __A14_2__IL03_n, S03_n, IL04, S04, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U14059(S04_n, __A14_2__IL04_n, S05, IL05, S05_n, __A14_2__IL05_n, GND, IL06, S06, __A14_2__IL06_n, S06_n, IL07, S07, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U14060(CLROPE, MYCLMP, __A14_NET_211,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15001(__A15_NET_200, WL16_n, WFBG_n, __A15_1__FB16, __A15_1__FB16_n, CFBG, GND, __A15_1__FB16_n, RFBG_n, __A15_1__BK16, WL14_n, WFBG_n, __A15_NET_198, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U15002(__A15_NET_200, __A15_NET_201, SUMA16_n, U2BBKG_n, SUMB16_n, __A15_NET_201, GND, __A15_NET_199, SUMA14_n, U2BBKG_n, SUMB14_n, __A15_1__FB16_n, __A15_1__FB16, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15003(__A15_1__BK16, __A15_NET_195, __A15_1__BK16, __A15_NET_197, __A15_NET_206, __A15_NET_207, GND, __A15_NET_202, __A15_NET_204, __A15_NET_192, __A15_NET_165, __A15_NET_210, __A15_NET_149, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U15004(__A15_NET_195, RL16_n_U15004_2, __A15_NET_197, RL15_n_U15004_4, __A15_NET_207, RL14_n_U15004_6, GND, RL13_n_U15004_8, __A15_NET_202, RL12_n_U15004_10, __A15_NET_189, RL11_n_U15004_12, __A15_NET_188, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b1) U15005(__A15_NET_198, __A15_NET_199, SUMA13_n, U2BBKG_n, SUMB13_n, __A15_NET_209, GND, __A15_1__FB13_n, __A15_NET_208, __A15_NET_209, __A15_1__FB13, __A15_1__FB14_n, __A15_1__FB14, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15006(__A15_1__FB14, __A15_1__FB14_n, CFBG, __A15_NET_206, __A15_1__FB14_n, RFBG_n, GND, WL13_n, WFBG_n, __A15_NET_208, __A15_1__FB13_n, CFBG, __A15_1__FB13, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15007(__A15_NET_204, __A15_1__FB13_n, RFBG_n, __A15_NET_203, WL12_n, WFBG_n, GND, __A15_1__FB12_n, CFBG, __A15_1__FB12, __A15_1__FB12_n, RFBG_n, __A15_NET_161, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U15008(SUMA12_n, U2BBKG_n, __A15_NET_203, __A15_NET_205, __A15_1__FB12, __A15_1__FB12_n, GND, __A15_NET_189, RSTRT, __A15_NET_161, __A15_1__RPTA12, __A15_NET_205, SUMB12_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15009(__A15_NET_162, WFBG_n, WL11_n, __A15_1__FB11, __A15_1__FB11_n, CFBG, GND, __A15_1__FB11_n, RFBG_n, __A15_NET_157, __A15_NET_157, __A15_NET_166, __A15_NET_188, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U15010(SUMA11_n, U2BBKG_n, __A15_NET_162, __A15_NET_163, __A15_1__FB11, __A15_1__FB11_n, GND, __A15_NET_158, SUMA03_n, U2BBKG_n, SUMB03_n, __A15_NET_163, SUMB11_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15011(__A15_NET_159, WL11_n, WEBG_n, __A15_NET_160, WL03_n, WBBEG_n, GND, EB11_n, CEBG, __A15_1__EB11, REBG_n, EB11_n, __A15_NET_166, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U15012(EB11_n, __A15_NET_158, __A15_NET_159, __A15_NET_160, __A15_1__EB11,  , GND,  , __A15_NET_167, __A15_NET_168, __A15_NET_164, EB10, __A15_1__EB10_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15013(__A15_1__BBK3, EB11_n, RBBEG_n, __A15_NET_168, WL10_n, WEBG_n, GND, WL02_n, WBBEG_n, __A15_NET_164, __A15_1__EB10_n, CEBG, EB10, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15014(SUMA02_n, U2BBKG_n, SUMA01_n, U2BBKG_n, SUMB01_n, __A15_NET_150, GND, __A15_1__F14, __A15_NET_153, __A15_NET_154, __A15_1__FB14_n, __A15_NET_167, SUMB02_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15015(__A15_NET_165, REBG_n, __A15_1__EB10_n, __A15_1__BBK2, __A15_1__EB10_n, RBBEG_n, GND, WL09_n, WEBG_n, __A15_NET_151, WL01_n, WBBEG_n, __A15_NET_152, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U15016(__A15_NET_192, RL10_n_U15016_2, __A15_NET_210, RL09_n_U15016_4, __A15_NET_181, RL06_n_U15016_6, GND, __A15_NET_229_U15016_8, __A15_NET_294, __A15_NET_229_U15016_10, __A15_NET_296, __A15_NET_232_U15016_12, __A15_NET_291, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U15017(__A15_1__EB9_n, __A15_NET_150, __A15_NET_151, __A15_NET_152, EB9,  , GND,  , __A15_1__FB14_n, __A15_1__FB16_n, E7_n, __A15_NET_153, __A15_1__F16, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15018(EB9, __A15_1__EB9_n, CEBG, __A15_NET_149, REBG_n, __A15_1__EB9_n, GND, __A15_1__EB9_n, RBBEG_n, __A15_1__BBK1, __A15_1__FB11_n, __A15_NET_153, __A15_NET_155, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15019(S12_n, __A15_NET_153, __A15_1__F11_n, __A15_1__F11, __A15_1__F12_n, __A15_1__F12, GND, __A15_1__F13_n, __A15_1__F13, __A15_1__F14_n, __A15_1__F14, __A15_1__F15_n, __A15_1__F15, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15020(__A15_1__F11_n, __A15_NET_155, __A15_NET_156, __A15_NET_156, S11_n, S12_n, GND, __A15_NET_153, __A15_1__FB12, __A15_1__F12_n, __A15_NET_153, __A15_1__FB13_n, __A15_1__F13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15021(E5, __A15_1__FB16_n, __A15_1__FB16_n, __A15_NET_184, __A15_NET_153, __A15_1__F15, GND, __A15_NET_184, E7_n, __A15_1__FB14_n, E6, __A15_NET_154, E7_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15022(__A15_1__F16, __A15_1__F16_n, __A15_NET_305, __A15_NET_301, KRPT, __A15_1__KRPTA_n, GND, __A15_NET_245, __A15_NET_244, __A15_NET_213, __A15_NET_224, __A15_1__PRPOR1, __A15_NET_218, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15023(XB4_n, XT4_n, __A15_1__KRPTA_n, XB0_n, XT5_n, __A15_NET_186, GND, __A15_NET_175, __A15_NET_185, __A15_NET_187, GOJAM, __A15_NET_187, __A15_1__KRPTA_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0) U15024(__A15_NET_185, RADRPT, __A15_NET_175, __A15_NET_174, HNDRPT, __A15_NET_171, GND, __A15_NET_179, __A15_1__RRPA1_n, __A15_1__RPTAD6, __A15_1__RRPA1_n, __A15_NET_177, __A15_1__RPTA12, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15025(__A15_NET_174, __A15_NET_186, __A15_1__PRPOR1, __A15_NET_185, __A15_1__DNRPTA, __A15_1__PRPOR3, GND, __A15_NET_179, __A15_1__PRPOR2, __A15_1__PRPOR3, __A15_1__PRPOR4, __A15_NET_171, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U15026(__A15_1__PRPOR4, __A15_1__PRPOR1, __A15_1__DNRPTA, __A15_NET_175, __A15_NET_174,  , GND,  , __A15_NET_171, __A15_NET_175, __A15_1__PRPOR1, __A15_1__DNRPTA, __A15_NET_177, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U15027(__A15_NET_181, CAD6, __A15_1__RPTAD6, __A15_NET_176, __A15_NET_177, RUPTOR_n, GND, __A15_NET_176, T10, RUPTOR_n, WOVR_n, OVF_n, __A15_NET_305, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15028(CA3_n, XB1_n, __A15_NET_306, GOJAM, __A15_NET_307, __A15_NET_295, GND, __A15_NET_307, XT0_n, XB4_n, __A15_1__KRPTA_n, T6RPT, ZOUT_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b1) U15029(__A15_NET_306, T6RPT, __A15_NET_295, __A15_NET_238, __A15_NET_302, __A15_NET_240, GND, __A15_NET_303, __A15_NET_243, __A15_NET_239, __A15_NET_236, __A15_NET_223, __A15_NET_237, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15030(CA3_n, XB0_n, __A15_NET_238, GOJAM, __A15_NET_300, __A15_NET_240, GND, __A15_NET_300, XB0_n, XT1_n, __A15_1__KRPTA_n, __A15_NET_302, __A15_NET_301, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15031(CA2_n, XB6_n, __A15_NET_239, GOJAM, __A15_NET_304, __A15_NET_243, GND, __A15_NET_304, XT1_n, XB4_n, __A15_1__KRPTA_n, __A15_NET_303, __A15_NET_301, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15032(CA2_n, XB7_n, __A15_NET_237, GOJAM, __A15_NET_235, __A15_NET_223, GND, __A15_NET_235, XT2_n, XB0_n, __A15_1__KRPTA_n, __A15_NET_236, __A15_NET_301, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b1, 1'b0) U15033(__A15_NET_234, KYRPT1, __A15_NET_225, __A15_NET_215, UPRUPT, __A15_NET_219, GND, DLKPLS, __A15_1__DNRPTA, __A15_NET_220, __A15_NET_295, __A15_NET_238, __A15_NET_241, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U15034(__A15_NET_234, GOJAM, XB4_n, XT2_n, __A15_1__KRPTA_n, __A15_2__KY1RST, GND, __A15_NET_226, KYRPT2, MKRPT, __A15_NET_217, __A15_NET_225, __A15_2__KY1RST, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15035(__A15_NET_226, GOJAM, XT3_n, XB0_n, __A15_1__KRPTA_n, __A15_2__KY2RST, GND, __A15_NET_219, __A15_NET_215, GOJAM, __A15_NET_246, __A15_NET_217, __A15_2__KY2RST, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15036(XT3_n, XB4_n, __A15_NET_220, GOJAM, DRPRST, __A15_1__DNRPTA, GND, DRPRST, XB0_n, XT4_n, __A15_1__KRPTA_n, __A15_NET_246, __A15_1__KRPTA_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15037(__A15_NET_294, __A15_NET_295, __A15_NET_242, __A15_NET_291, __A15_NET_241, __A15_NET_242, GND, __A15_NET_245, __A15_NET_237, __A15_NET_222, __A15_NET_213, __A15_NET_226, __A15_NET_216, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15038(__A15_NET_221, __A15_NET_214, __A15_NET_295, __A15_NET_239, __A15_NET_240, __A15_NET_242, GND, __A15_NET_290, __A15_NET_216, __A15_NET_214, __A15_1__PRPOR4, __A15_NET_296, __A15_1__PRPOR3, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U15039(__A15_NET_290, __A15_NET_232_U15039_2, __A15_NET_265, RL03_n_U15039_4, __A15_NET_297, RL04_n_U15039_6, GND, RL05_n_U15039_8, __A15_NET_298, RL02_n_U15039_10, __A15_NET_299, RL01_n_U15039_12, __A15_NET_310, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15040(__A15_NET_295, __A15_NET_243, __A15_NET_245, __A15_NET_234, __A15_NET_223, __A15_NET_221, GND, __A15_NET_224, __A15_NET_245, __A15_NET_225, __A15_NET_223, __A15_NET_244, __A15_NET_240, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U15041(__A15_NET_260, __A15_NET_221, __A15_NET_222, __A15_NET_216, __A15_NET_214,  , GND,  , __A15_2__RPTAD3, __A15_1__BBK3, CAD3, R6, __A15_NET_265, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15042(__A15_NET_213, __A15_NET_215, __A15_NET_213, __A15_NET_219, __A15_NET_217, __A15_NET_218, GND,  ,  ,  ,  , __A15_NET_214, __A15_NET_217, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15043(__A15_1__PRPOR2, __A15_1__PRPOR1, __A15_NET_220, __A15_2__RPTAD3, __A15_1__RRPA1_n, __A15_NET_229, GND, __A15_1__RRPA1_n, __A15_NET_232, __A15_2__RPTAD4, __A15_2__RPTAD4, CAD4, __A15_NET_297, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15044(RRPA, __A15_1__RRPA1_n, STRGAT, __A15_NET_227, __A15_1__F11, __A15_NET_228, GND, __A15_NET_272, __A15_1__F11_n, __A15_NET_273, S10, __A15_NET_271, S10_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15045(__A15_NET_298, __A15_2__RPTAD5, CAD5, __A15_2__RPTAD5, __A15_1__RRPA1_n, __A15_NET_260, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15046(CAD2, __A15_1__BBK2, CAD1, __A15_1__BBK1, RB1F, __A15_NET_310, GND, STR412, __A15_NET_227, __A15_NET_273, __A15_NET_228, __A15_NET_299, R6, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15047(__A15_NET_227, __A15_NET_271, __A15_NET_227, __A15_NET_273, __A15_NET_272, STR210, GND, STR19, __A15_NET_227, __A15_NET_271, __A15_NET_272, STR311, __A15_NET_228, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15048(__A15_NET_274, __A15_1__F16, __A15_1__F15, __A15_NET_269, __A15_1__F16, __A15_1__F15_n, GND, __A15_1__F15, __A15_1__F16_n, __A15_NET_287, __A15_2__NE036_n, __A15_1__F12, __A15_2__036L, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15049(__A15_NET_274, __A15_NET_268, __A15_1__F14_n, __A15_NET_270, __A15_1__F13_n, __A15_NET_285, GND, __A15_NET_282, __A15_1__F13, __A15_NET_284, __A15_1__F14, __A15_NET_283, __A15_NET_269, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15050(__A15_NET_268, __A15_NET_270, __A15_NET_268, __A15_NET_270, __A15_NET_282, __A15_2__NE01, GND, __A15_2__NE02, __A15_NET_268, __A15_NET_284, __A15_NET_285, __A15_2__NE00, __A15_NET_285, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15051(__A15_NET_268, __A15_NET_284, __A15_NET_283, __A15_NET_270, __A15_NET_285, __A15_2__NE04, GND, __A15_2__NE05, __A15_NET_283, __A15_NET_270, __A15_NET_282, __A15_2__NE03, __A15_NET_282, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15052(__A15_NET_283, __A15_NET_284, __A15_NET_283, __A15_NET_284, __A15_NET_282, __A15_2__NE07, GND, __A15_2__NE10, __A15_NET_286, __A15_NET_270, __A15_NET_285, __A15_2__NE06, __A15_NET_285, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15053(__A15_NET_287, __A15_NET_286, __A15_NET_251, STR14, __A15_2__NE012_n, ROPER, GND, LOMOD, __A15_NET_266, STR58, __A15_NET_267, ROPES, __A15_2__NE345_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15054(__A15_2__NE00, __A15_2__NE03, __A15_2__NE00, __A15_2__NE01, __A15_2__NE02, __A15_2__NE012_n, GND, __A15_2__NE147_n, __A15_2__NE01, __A15_2__NE04, __A15_2__NE07, __A15_2__NE036_n, __A15_2__NE06, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15055(__A15_2__NE04, __A15_2__NE03, __A15_2__NE02, __A15_2__NE05, __A15_2__NE10, __A15_2__NE2510_n, GND, __A15_2__NE6710_n, __A15_2__NE06, __A15_2__NE07, __A15_2__NE10, __A15_2__NE345_n, __A15_2__NE05, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15056(__A15_2__147H, __A15_2__NE147_n, __A15_1__F12_n, __A15_2__2510L, __A15_2__NE2510_n, __A15_1__F12, GND, __A15_2__NE036_n, __A15_1__F12_n, __A15_2__036H, __A15_2__NE147_n, __A15_1__F12, __A15_2__147L, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U15057(__A15_2__2510H, __A15_2__NE2510_n, __A15_1__F12_n, __A15_NET_251, __A15_2__036L, __A15_2__147H, GND, __A15_2__2510L, __A15_2__036H, __A15_NET_267, __A15_2__147L, __A15_2__2510H, __A15_NET_262, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U15058(__A15_2__036L, __A15_2__147L, __A15_2__147H, __A15_2__2510H, __A15_2__2510L, __A15_NET_261, GND,  ,  ,  ,  , __A15_NET_266, __A15_2__036H, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U15059(__A15_NET_261, HIMOD, __A15_NET_262, STR912, __A15_2__NE6710_n, ROPET, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16001(__A16_NET_181, CHWL01_n, __A16_1__WCH05_n, __A16_NET_191, __A16_NET_181, __A16_NET_182, GND, __A16_NET_191, __A16_1__CCH05, __A16_NET_182, __A16_NET_191, __A16_1__RCH05_n, __A16_NET_183, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16002(__A16_NET_191, __A16_1__RCpXpP, __A16_NET_175, __A16_1__RCpZpR, __A16_NET_180, __A16_1__RCmXmP, GND, __A16_1__RCmZmR, __A16_NET_127, __A16_1__RCmXpP, __A16_NET_126, __A16_1__RCmZpR, __A16_NET_136, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16003(__A16_NET_177, __A16_NET_183, __A16_NET_128, __A16_NET_123, CH3202, __A16_NET_187, GND, __A16_NET_186, __A16_NET_137, __A16_NET_133, CH3203, __A16_NET_184, CH3201, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U16004(__A16_NET_184, CHOR01_n_U16004_2, __A16_NET_187, CHOR02_n_U16004_4, __A16_NET_186, CHOR03_n_U16004_6, GND, CHOR04_n_U16004_8, __A16_NET_172, CHOR05_n_U16004_10, __A16_NET_174, CHOR06_n_U16004_12, __A16_NET_173, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16005(__A16_NET_185, CHWL01_n, __A16_1__WCH06_n, __A16_NET_175, __A16_NET_185, __A16_NET_176, GND, __A16_NET_175, __A16_1__CCH06, __A16_NET_176, __A16_NET_175, __A16_1__RCH06_n, __A16_NET_177, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16006(__A16_NET_178, CHWL02_n, __A16_1__WCH05_n, __A16_NET_180, __A16_NET_178, __A16_NET_179, GND, __A16_NET_180, __A16_1__CCH05, __A16_NET_179, __A16_NET_180, __A16_1__RCH05_n, __A16_NET_123, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16007(__A16_NET_124, CHWL02_n, __A16_1__WCH06_n, __A16_NET_127, __A16_NET_124, __A16_NET_125, GND, __A16_NET_127, __A16_1__CCH06, __A16_NET_125, __A16_NET_127, __A16_1__RCH06_n, __A16_NET_128, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16008(__A16_NET_121, CHWL03_n, __A16_1__WCH05_n, __A16_NET_126, __A16_NET_121, __A16_NET_122, GND, __A16_NET_126, __A16_1__CCH05, __A16_NET_122, __A16_NET_126, __A16_1__RCH05_n, __A16_NET_133, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16009(__A16_NET_134, CHWL03_n, __A16_1__WCH06_n, __A16_NET_136, __A16_NET_134, __A16_NET_135, GND, __A16_NET_136, __A16_1__CCH06, __A16_NET_135, __A16_NET_136, __A16_1__RCH06_n, __A16_NET_137, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16010(__A16_NET_130, CHWL04_n, __A16_1__WCH05_n, __A16_NET_131, __A16_NET_130, __A16_NET_129, GND, __A16_NET_131, __A16_1__CCH05, __A16_NET_129, __A16_NET_131, __A16_1__RCH05_n, __A16_NET_132, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16011(__A16_NET_131, __A16_1__RCpXmP, __A16_NET_111, __A16_1__RCpZmR, __A16_NET_104, __A16_1__RCpXpY, GND, __A16_1__RCpYpR, __A16_NET_120, __A16_1__RCmXmY, __A16_NET_115, __A16_1__RCmYmR, __A16_NET_159, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16012(__A16_NET_112, __A16_NET_132, __A16_NET_119, __A16_NET_105, CH3205, __A16_NET_174, GND, __A16_NET_173, __A16_NET_160, __A16_NET_116, CH3206, __A16_NET_172, CH3204, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16013(__A16_NET_108, CHWL04_n, __A16_1__WCH06_n, __A16_NET_111, __A16_NET_108, __A16_NET_109, GND, __A16_NET_111, __A16_1__CCH06, __A16_NET_109, __A16_NET_111, __A16_1__RCH06_n, __A16_NET_112, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16014(__A16_NET_103, CHWL05_n, __A16_1__WCH05_n, __A16_NET_104, __A16_NET_103, __A16_NET_102, GND, __A16_NET_104, __A16_1__CCH05, __A16_NET_102, __A16_NET_104, __A16_1__RCH05_n, __A16_NET_105, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16015(__A16_NET_106, CHWL05_n, __A16_1__WCH06_n, __A16_NET_120, __A16_NET_106, __A16_NET_107, GND, __A16_NET_120, __A16_1__CCH06, __A16_NET_107, __A16_NET_120, __A16_1__RCH06_n, __A16_NET_119, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16016(__A16_NET_113, CHWL06_n, __A16_1__WCH05_n, __A16_NET_115, __A16_NET_113, __A16_NET_114, GND, __A16_NET_115, __A16_1__CCH05, __A16_NET_114, __A16_NET_115, __A16_1__RCH05_n, __A16_NET_116, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16017(__A16_NET_117, CHWL06_n, __A16_1__WCH06_n, __A16_NET_159, __A16_NET_117, __A16_NET_118, GND, __A16_NET_159, __A16_1__CCH06, __A16_NET_118, __A16_NET_159, __A16_1__RCH06_n, __A16_NET_160, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16018(__A16_NET_163, CHWL07_n, __A16_1__WCH05_n, __A16_NET_154, __A16_NET_163, __A16_NET_153, GND, __A16_NET_154, __A16_1__CCH05, __A16_NET_153, __A16_NET_154, __A16_1__RCH05_n, __A16_NET_155, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16019(__A16_NET_154, __A16_1__RCmXpY, __A16_NET_157, __A16_1__RCmYpR, __A16_NET_164, __A16_1__RCpXmY, GND, __A16_1__RCpYmR, __A16_NET_168, __A16_1__WCH05_n, __A16_NET_144, __A16_1__WCH06_n, __A16_NET_145, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16020(__A16_NET_169, __A16_NET_155, __A16_NET_143, __A16_NET_165, CH3208, __A16_NET_193, GND, __A16_NET_144, WCHG_n, XT0_n, XB5_n, __A16_NET_192, CH3207, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U16021(__A16_NET_192, CHOR07_n_U16021_2, __A16_NET_193, CHOR08_n_U16021_4, __A16_NET_249, CHOR01_n_U16021_6, GND, CHOR02_n_U16021_8, __A16_NET_268, CHOR03_n_U16021_10, __A16_NET_243, CHOR04_n_U16021_12, __A16_NET_242, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16022(__A16_NET_152, CHWL07_n, __A16_1__WCH06_n, __A16_NET_157, __A16_NET_152, __A16_NET_156, GND, __A16_NET_157, __A16_1__CCH06, __A16_NET_156, __A16_NET_157, __A16_1__RCH06_n, __A16_NET_169, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16023(__A16_NET_170, CHWL08_n, __A16_1__WCH05_n, __A16_NET_164, __A16_NET_170, __A16_NET_171, GND, __A16_NET_164, __A16_1__CCH05, __A16_NET_171, __A16_NET_164, __A16_1__RCH05_n, __A16_NET_165, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16024(__A16_NET_166, CHWL08_n, __A16_1__WCH06_n, __A16_NET_168, __A16_NET_166, __A16_NET_167, GND, __A16_NET_168, __A16_1__CCH06, __A16_NET_167, __A16_NET_168, __A16_1__RCH06_n, __A16_NET_143, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16025(WCHG_n, XT0_n, CCHG_n, XT0_n, XB5_n, __A16_NET_138, GND, __A16_NET_140, CCHG_n, XT0_n, XB6_n, __A16_NET_145, XB6_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16026(__A16_NET_110, __A16_1__CCH05, __A16_NET_139, __A16_1__RCH05_n, __A16_NET_142, __A16_1__RCH06_n, GND, __A16_1__CCH06, __A16_NET_141, __A16_1__TVCNAB, __A16_NET_150, __A16_1__OT1207, __A16_NET_146, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U16027(__A16_NET_110, __A16_NET_138, GOJAM, __A16_NET_139, XT0_n, XB5_n, GND, XT0_n, XB6_n, __A16_NET_142, __A16_NET_140, GOJAM, __A16_NET_141, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16028(__A16_NET_148, CHWL08_n, WCH12_n, __A16_NET_150, __A16_NET_148, __A16_NET_149, GND, __A16_NET_150, CCH12, __A16_NET_149, RCH12_n, __A16_NET_150, CH1208, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16029(__A16_NET_151, WCH12_n, CHWL07_n, __A16_NET_146, __A16_NET_151, __A16_NET_147, GND, __A16_NET_146, CCH12, __A16_NET_147, RCH12_n, __A16_NET_146, __A16_1__CH1207, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16030(__A16_NET_147, __A16_1__OT1207_n, __A16_NET_274, __A16_2__ZOPCDU, __A16_NET_273, __A16_2__ISSWAR, GND, __A16_2__ENEROP, __A16_NET_252, COMACT, __A16_NET_270, __A16_2__STARON, __A16_NET_271, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16031(__A16_NET_255, CHWL01_n, WCH12_n, __A16_NET_274, __A16_NET_255, __A16_NET_256, GND, __A16_NET_274, CCH12, __A16_NET_256, __A16_NET_274, RCH12_n, __A16_NET_257, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16032(__A16_NET_257, __A16_NET_250, __A16_NET_254, __A16_NET_267, CH1502, __A16_NET_268, GND, __A16_NET_243, __A16_NET_261, __A16_NET_264, CH1503, __A16_NET_249, CH1501, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16033(__A16_NET_258, CHWL01_n, WCH11_n, __A16_NET_273, __A16_NET_258, __A16_NET_259, GND, __A16_NET_273, CCH11, __A16_NET_259, __A16_NET_273, RCH11_n, __A16_NET_250, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16034(__A16_NET_251, CHWL02_n, WCH12_n, __A16_NET_252, __A16_NET_251, __A16_NET_253, GND, __A16_NET_252, CCH12, __A16_NET_253, __A16_NET_252, RCH12_n, __A16_NET_254, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16035(__A16_NET_265, CHWL02_n, WCH11_n, __A16_NET_270, __A16_NET_265, __A16_NET_266, GND, __A16_NET_270, CCH11, __A16_NET_266, __A16_NET_270, RCH11_n, __A16_NET_267, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16036(__A16_NET_269, CHWL03_n, WCH12_n, __A16_NET_271, __A16_NET_269, __A16_NET_260, GND, __A16_NET_271, CCH12, __A16_NET_260, __A16_NET_271, RCH12_n, __A16_NET_261, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16037(__A16_NET_262, CHWL03_n, WCH11_n, __A16_NET_272, __A16_NET_262, __A16_NET_263, GND, __A16_NET_272, CCH11, __A16_NET_263, __A16_NET_272, RCH11_n, __A16_NET_264, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16038(__A16_NET_272, UPLACT, __A16_NET_246, __A16_2__COARSE, __A16_NET_212, TMPOUT, GND, __A16_2__ZIMCDU, __A16_NET_211, __A16_2__ENERIM, __A16_NET_220, __A16_2__S4BTAK, __A16_NET_197, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16039(__A16_NET_244, CHWL04_n, WCH12_n, __A16_NET_246, __A16_NET_244, __A16_NET_245, GND, __A16_NET_246, CCH12, __A16_NET_245, __A16_NET_246, RCH12_n, __A16_NET_216, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16040(__A16_NET_213, CHWL04_n, WCH11_n, __A16_NET_212, __A16_NET_213, __A16_NET_214, GND, __A16_NET_212, CCH11, __A16_NET_214, __A16_NET_212, RCH11_n, __A16_NET_217, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16041(__A16_NET_216, __A16_NET_217, __A16_NET_225, __A16_NET_226, CH0705, __A16_NET_248, GND, __A16_NET_247, __A16_NET_198, __A16_NET_199, CH0706, __A16_NET_242, CH1504, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16042(__A16_NET_209, CHWL05_n, WCH12_n, __A16_NET_211, __A16_NET_209, __A16_NET_210, GND, __A16_NET_211, CCH12, __A16_NET_210, __A16_NET_211, RCH12_n, __A16_NET_225, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16043(__A16_NET_215, CHWL05_n, WCH11_n, __A16_NET_224, __A16_NET_215, __A16_NET_223, GND, __A16_NET_224, CCH11, __A16_NET_223, __A16_NET_224, RCH11_n, __A16_NET_226, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U16044(__A16_NET_248, CHOR05_n_U16044_2, __A16_NET_247, CHOR06_n_U16044_4, __A16_NET_238, CHOR07_n_U16044_6, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16045(__A16_NET_218, CHWL06_n, WCH12_n, __A16_NET_220, __A16_NET_218, __A16_NET_219, GND, __A16_NET_220, CCH12, __A16_NET_219, __A16_NET_220, RCH12_n, __A16_NET_198, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16046(__A16_NET_221, CHWL06_n, WCH11_n, __A16_NET_196, __A16_NET_221, __A16_NET_222, GND, __A16_NET_196, CCH11, __A16_NET_222, __A16_NET_196, RCH11_n, __A16_NET_199, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U16047(KYRLS, __A16_NET_224, FLASH, VNFLSH, __A16_NET_196, FLASH_n, GND, __A16_NET_235, FLASH, OPEROR, __A16_NET_229, GOJAM, __A16_NET_233, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16048(__A16_NET_195, CHWL09_n, WCH12_n, __A16_NET_197, __A16_NET_195, __A16_NET_194, GND, __A16_NET_197, CCH12, __A16_NET_194, __A16_NET_197, RCH12_n, CH1209, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16049(__A16_NET_206, CHWL10_n, WCH12_n, __A16_NET_205, __A16_NET_206, __A16_NET_204, GND, __A16_NET_205, CCH12, __A16_NET_204, __A16_NET_205, RCH12_n, CH1210, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16050(__A16_NET_205, __A16_2__ZEROPT, __A16_NET_200, __A16_2__DISDAC, __A16_NET_240, __A16_2__MROLGT, GND, __A16_2__S4BSEQ, __A16_NET_228, __A16_2__S4BOFF, __A16_NET_232, WCH12_n, __A16_NET_227, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16051(__A16_NET_207, CHWL11_n, WCH12_n, __A16_NET_200, __A16_NET_207, __A16_NET_208, GND, __A16_NET_200, CCH12, __A16_NET_208, __A16_NET_200, RCH12_n, CH1211, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16052(__A16_NET_201, CHWL07_n, WCH11_n, __A16_NET_235, __A16_NET_201, __A16_NET_202, GND, __A16_NET_235, CCH11, __A16_NET_202, __A16_NET_235, RCH11_n, __A16_NET_203, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U16053(__A16_1__CH1207, __A16_NET_203, WCHG_n, XB2_n, XT1_n, __A16_NET_227, GND, __A16_NET_229, CCHG_n, XB2_n, XT1_n, __A16_NET_238, CH0707, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16054(__A16_NET_236, CHWL12_n, WCH12_n, __A16_NET_240, __A16_NET_236, __A16_NET_237, GND, __A16_NET_240, CCH12, __A16_NET_237, __A16_NET_240, RCH12_n, CH1212, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16055(__A16_NET_239, CHWL13_n, WCH12_n, __A16_NET_228, __A16_NET_239, __A16_NET_241, GND, __A16_NET_228, CCH12, __A16_NET_241, __A16_NET_228, RCH12_n, CH1213, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U16056(__A16_NET_230, CHWL14_n, WCH12_n, __A16_NET_232, __A16_NET_230, __A16_NET_231, GND, __A16_NET_232, CCH12, __A16_NET_231, __A16_NET_232, RCH12_n, CH1214, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U16057(__A16_NET_233, CCH12, __A16_NET_234, RCH12_n,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U16058(__A16_NET_234, XT1_n, XB2_n,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17001(__A17_NET_250, IN3301, RCH33_n, __A17_NET_249, XB3_n, XT3_n, GND, ULLTHR, __A17_1__RCH30_n, __A17_NET_248, XB0_n, XT3_n, __A17_NET_215, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U17002(__A17_NET_249, RCH33_n, __A17_NET_215, __A17_1__RCH30_n, __A17_NET_251, __A17_1__RCH31_n, GND, __A17_1__RCH32_n, __A17_NET_204, __A17_1__F04B_n, F04B, RLYB01, __A17_NET_329, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17003(__A17_NET_246, CHOR01_n_U17003_2, __A17_NET_238, CHOR02_n_U17003_4, __A17_NET_242, CHOR03_n_U17003_6, GND, CHOR04_n_U17003_8, __A17_NET_258, CHOR05_n_U17003_10, __A17_NET_256, CHOR06_n_U17003_12, __A17_NET_253, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17004(__A17_NET_247, MANpP, __A17_1__RCH31_n, __A17_NET_251, XB1_n, XT3_n, GND, SMSEPR, __A17_1__RCH30_n, __A17_NET_240, RRPONA, RCH33_n, __A17_NET_241, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17005(__A17_NET_239, MANmP, __A17_1__RCH31_n, __A17_NET_245, RRRLSC, RCH33_n, GND, MANpY, __A17_1__RCH31_n, __A17_NET_243, SPSRDY, __A17_1__RCH30_n, __A17_NET_244, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17006(__A17_NET_250, __A17_NET_248, __A17_NET_241, __A17_NET_240, __A17_NET_239, __A17_NET_238, GND, __A17_NET_242, __A17_NET_245, __A17_NET_244, __A17_NET_243, __A17_NET_246, __A17_NET_247, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17007(__A17_NET_263, S4BSAB, __A17_1__RCH30_n, __A17_NET_260, ZEROP, RCH33_n, GND, MANmY, __A17_1__RCH31_n, __A17_NET_259, LFTOFF, __A17_1__RCH30_n, __A17_NET_261, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17008(__A17_NET_260, __A17_NET_263, __A17_NET_262, __A17_NET_261, __A17_NET_264, __A17_NET_256, GND, __A17_NET_253, __A17_NET_254, __A17_NET_252, __A17_NET_255, __A17_NET_258, __A17_NET_259, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17009(__A17_NET_262, OPMSW2, RCH33_n, __A17_NET_264, MANpR, __A17_1__RCH31_n, GND, GUIREL, __A17_1__RCH30_n, __A17_NET_252, OPMSW3, RCH33_n, __A17_NET_254, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17010(__A17_NET_255, MANmR, __A17_1__RCH31_n, __A17_NET_237, OPCDFL, __A17_1__RCH30_n, GND, STRPRS, RCH33_n, __A17_NET_257, TRANpX, __A17_1__RCH31_n, __A17_NET_229, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17011(__A17_NET_257, __A17_NET_237, __A17_NET_227, __A17_NET_232, __A17_NET_231, __A17_NET_230, GND, __A17_NET_225, __A17_NET_198, __A17_NET_197, __A17_NET_196, __A17_NET_228, __A17_NET_229, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17012(__A17_NET_228, CHOR07_n_U17012_2, __A17_NET_230, CHOR08_n_U17012_4, __A17_NET_225, CHOR09_n_U17012_6, GND, CHOR10_n_U17012_8, __A17_NET_226, CHOR11_n_U17012_10, __A17_NET_235, CHOR12_n_U17012_12, __A17_NET_236, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17013(__A17_NET_232, IN3008, __A17_1__RCH30_n, __A17_NET_227, LVDAGD, RCH33_n, GND, TRANmX, __A17_1__RCH31_n, __A17_NET_231, IMUOPR, __A17_1__RCH30_n, __A17_NET_197, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17014(__A17_NET_198, LRRLSC, RCH33_n, __A17_NET_196, TRANpY, __A17_1__RCH31_n, GND, CTLSAT, __A17_1__RCH30_n, __A17_NET_200, TRANmY, __A17_1__RCH31_n, __A17_NET_199, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17015(CH3310, __A17_NET_200, __A17_NET_192, __A17_NET_191, __A17_NET_190, __A17_NET_235, GND, __A17_NET_236, __A17_NET_195, __A17_NET_193, __A17_NET_194, __A17_NET_226, __A17_NET_199, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17016(__A17_NET_191, IMUCAG, __A17_1__RCH30_n, __A17_NET_192, LEMATT, __A17_1__RCH32_n, GND, TRANpZ, __A17_1__RCH31_n, __A17_NET_190, CDUFAL, __A17_1__RCH30_n, __A17_NET_193, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17017(__A17_NET_195, IN3212, __A17_1__RCH32_n, __A17_NET_194, TRANmZ, __A17_1__RCH31_n, GND, IMUFAL, __A17_1__RCH30_n, __A17_NET_207, IN3213, __A17_1__RCH32_n, __A17_NET_208, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17018(__A17_NET_208, __A17_NET_207, __A17_NET_210, __A17_NET_209, __A17_NET_203, __A17_NET_234, GND, __A17_NET_267, __A17_NET_202, __A17_NET_201, __A17_NET_205, __A17_NET_233, __A17_NET_206, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17019(__A17_NET_233, CHOR13_n_U17019_2, __A17_NET_234, CHOR14_n_U17019_4, __A17_NET_267, CHOR16_n_U17019_6, GND, __A17_NET_176_U17019_8, __A17_NET_266, __A17_NET_176_U17019_10, __A17_NET_265, __A17_NET_183_U17019_12, __A17_NET_270, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17020(__A17_NET_206, HOLFUN, __A17_1__RCH31_n, __A17_NET_209, ISSTOR, __A17_1__RCH30_n, GND, IN3214, __A17_1__RCH32_n, __A17_NET_210, FREFUN, __A17_1__RCH31_n, __A17_NET_203, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17021(__A17_NET_201, TEMPIN, __A17_1__RCH30_n, __A17_NET_202, IN3216, __A17_1__RCH32_n, GND, GCAPCL, __A17_1__RCH31_n, __A17_NET_205, XB2_n, XT3_n, __A17_NET_204, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17022(MANpP, MANmP, MANmY, MANpR, MANmR, __A17_NET_265, GND, __A17_NET_179, __A17_NET_180, __A17_NET_176, F05A_n, __A17_NET_266, MANpY, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U17023(__A17_NET_182, CHWL12_n, WCH13_n, __A17_NET_180, __A17_NET_182, __A17_NET_181, GND, __A17_NET_179, __A17_NET_178, __A17_NET_177, __A17_1__F04B_n, FS05_n, __A17_1__FO5D, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17024(__A17_NET_180, GOJAM, __A17_NET_177, __A17_NET_176, __A17_1__FO5D, __A17_NET_178, GND, __A17_NET_270, TRANpX, TRANmX, TRANpY, __A17_NET_181, __A17_1__TRP31A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U17025(__A17_1__TRP31A, __A17_NET_177, F05B_n, __A17_NET_185, __A17_NET_184, __A17_NET_186, GND, CHWL13_n, WCH13_n, __A17_NET_189, __A17_NET_185, F05B_n, __A17_1__TRP31B, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17026(TRANmY, TRANpZ, __A17_NET_187, __A17_NET_183, F05A_n, __A17_NET_184, GND, __A17_NET_186, __A17_NET_185, __A17_NET_183, __A17_1__FO5D, __A17_NET_269, TRANmZ, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17027(__A17_NET_269, __A17_NET_183_U17027_2, __A17_NET_217, __A17_NET_220_U17027_4, __A17_NET_222, __A17_NET_220_U17027_6, GND, __A17_NET_220_U17027_8, __A17_NET_221, CHOR01_n_U17027_10, __A17_NET_323, CHOR07_n_U17027_12, __A17_NET_338, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17028(__A17_NET_187, GOJAM, MNIMpR, MNIMmR, TRST9, __A17_NET_222, GND, __A17_NET_221, TRST10, PCHGOF, ROLGOF, __A17_NET_188, __A17_1__TRP31B, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17029(__A17_NET_187, __A17_NET_189, __A17_NET_188, CH3201, MNIMpP, __A17_1__RCH32_n, GND, MNIMmP, __A17_1__RCH32_n, CH3202, MNIMpY, __A17_1__RCH32_n, CH3203, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17030(CH3204, MNIMmY, __A17_1__RCH32_n, CH3205, MNIMpR, __A17_1__RCH32_n, GND, MNIMmR, __A17_1__RCH32_n, CH3206, TRST9, __A17_1__RCH32_n, CH3207, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U17031(CH3208, TRST10, __A17_1__RCH32_n, CH3209, PCHGOF, __A17_1__RCH32_n, GND, ROLGOF, __A17_1__RCH32_n, CH3210, __A17_NET_213, __A17_NET_212, __A17_NET_211, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U17032(__A17_NET_217, MNIMpP, MNIMmP, MNIMpY, MNIMmY,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17033(WCHG_n, XT1_n, __A17_NET_214, __A17_NET_220, F05A_n, __A17_NET_213, GND, __A17_NET_212, __A17_NET_211, __A17_1__FO5D, __A17_NET_220, __A17_NET_300, XB1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U17034(__A17_1__TRP32, __A17_NET_211, F05B_n, __A17_NET_219, CHWL14_n, WCH13_n, GND, __A17_NET_219, __A17_NET_218, __A17_NET_214, __A17_NET_216, TPOR_n, HNDRPT, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17035(__A17_NET_214, GOJAM, __A17_1__TRP31A, __A17_1__TRP31B, __A17_1__TRP32, __A17_NET_216, GND, __A17_NET_323, CH1301, __A17_NET_324, CH1401, __A17_NET_218, __A17_1__TRP32, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17036(CH3313, PIPAFL, RCH33_n, CH3314, AGCWAR, RCH33_n, GND, OSCALM, RCH33_n, CH3316, CHWL01_n, __A17_2__WCH10_n, __A17_NET_328, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17037(__A17_NET_329, __A17_NET_328, __A17_NET_327, __A17_NET_327, __A17_NET_329, __A17_2__CCH10, GND, __A17_NET_329, __A17_2__RCH10_n, __A17_NET_324, CHWL02_n, __A17_2__WCH10_n, __A17_NET_325, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17038(__A17_NET_332, __A17_NET_325, __A17_NET_326, __A17_NET_326, __A17_NET_332, __A17_2__CCH10, GND, __A17_NET_332, __A17_2__RCH10_n, __A17_NET_333, CHWL03_n, __A17_2__WCH10_n, __A17_NET_331, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U17039(__A17_NET_332, RLYB02, __A17_NET_314, RLYB03, __A17_NET_320, RLYB04, GND, RLYB05, __A17_NET_348, RLYB06, __A17_NET_355, RLYB07, __A17_NET_354, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17040(CH1302, __A17_NET_333, CH1303, __A17_NET_316, CH1403, __A17_NET_311, GND, __A17_NET_321, CH1304, __A17_NET_322, CH1404, __A17_NET_330, CH1402, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17041(__A17_NET_330, CHOR02_n_U17041_2, __A17_NET_311, CHOR03_n_U17041_4, __A17_NET_321, CHOR04_n_U17041_6, GND, CHOR05_n_U17041_8, __A17_NET_350, CHOR06_n_U17041_10, __A17_NET_356, CHOR08_n_U17041_12, __A17_NET_343, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17042(__A17_NET_314, __A17_NET_331, __A17_NET_315, __A17_NET_315, __A17_NET_314, __A17_2__CCH10, GND, __A17_NET_314, __A17_2__RCH10_n, __A17_NET_316, CHWL04_n, __A17_2__WCH10_n, __A17_NET_312, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17043(__A17_NET_320, __A17_NET_312, __A17_NET_313, __A17_NET_313, __A17_NET_320, __A17_2__CCH10, GND, __A17_NET_320, __A17_2__RCH10_n, __A17_NET_322, CHWL05_n, __A17_2__WCH10_n, __A17_NET_318, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17044(__A17_NET_348, __A17_NET_318, __A17_NET_319, __A17_NET_319, __A17_NET_348, __A17_2__CCH10, GND, __A17_NET_348, __A17_2__RCH10_n, __A17_NET_349, CHWL06_n, __A17_2__WCH10_n, __A17_NET_346, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17045(CH1305, __A17_NET_349, CH1306, __A17_NET_347, CH1406, __A17_NET_356, GND,  ,  ,  ,  , __A17_NET_350, CH1405, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17046(__A17_NET_355, __A17_NET_346, __A17_NET_344, __A17_NET_344, __A17_NET_355, __A17_2__CCH10, GND, __A17_NET_355, __A17_2__RCH10_n, __A17_NET_347, CHWL07_n, __A17_2__WCH10_n, __A17_NET_352, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17047(__A17_NET_354, __A17_NET_352, __A17_NET_351, __A17_NET_351, __A17_NET_354, __A17_2__CCH10, GND, __A17_NET_354, __A17_2__RCH10_n, __A17_NET_337, CHWL08_n, __A17_2__WCH10_n, __A17_NET_334, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17048(CH1307, __A17_NET_337, CH1308, __A17_NET_342, CH1408, __A17_NET_343, GND, __A17_NET_287, CH1309, __A17_NET_286, CH1409, __A17_NET_338, CH1407, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17049(__A17_NET_336, __A17_NET_334, __A17_NET_335, __A17_NET_335, __A17_NET_336, __A17_2__CCH10, GND, __A17_NET_336, __A17_2__RCH10_n, __A17_NET_342, CHWL09_n, __A17_2__WCH10_n, __A17_NET_339, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U17050(__A17_NET_336, RLYB08, __A17_NET_341, RLYB09, __A17_NET_283, RLYB10, GND, RLYB11, __A17_NET_289, RYWD12, __A17_NET_273, RYWD13, __A17_NET_281, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17051(__A17_NET_341, __A17_NET_339, __A17_NET_340, __A17_NET_340, __A17_NET_341, __A17_2__CCH10, GND, __A17_NET_341, __A17_2__RCH10_n, __A17_NET_286, CHWL10_n, __A17_2__WCH10_n, __A17_NET_288, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17052(__A17_NET_287, CHOR09_n_U17052_2, __A17_NET_285, CHOR10_n_U17052_4, __A17_NET_275, CHOR11_n_U17052_6, GND, CHOR12_n_U17052_8, __A17_NET_272, CHOR13_n_U17052_10, __A17_NET_278, CHOR14_n_U17052_12, __A17_NET_302, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17053(__A17_NET_283, __A17_NET_288, __A17_NET_282, __A17_NET_282, __A17_NET_283, __A17_2__CCH10, GND, __A17_NET_283, __A17_2__RCH10_n, __A17_NET_284, CHWL11_n, __A17_2__WCH10_n, __A17_NET_292, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17054(CH1310, __A17_NET_284, CH1311, __A17_NET_291, CH1411, __A17_NET_275, GND, __A17_NET_272, CH3312, __A17_NET_271, CH1412, __A17_NET_285, CH1410, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17055(__A17_NET_289, __A17_NET_292, __A17_NET_290, __A17_NET_290, __A17_NET_289, __A17_2__CCH10, GND, __A17_NET_289, __A17_2__RCH10_n, __A17_NET_291, CHWL12_n, __A17_2__WCH10_n, __A17_NET_276, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17056(__A17_NET_273, __A17_NET_276, __A17_NET_274, __A17_NET_274, __A17_NET_273, __A17_2__CCH10, GND, __A17_NET_273, __A17_2__RCH10_n, __A17_NET_271, CHWL13_n, __A17_2__WCH10_n, __A17_NET_279, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17057(__A17_NET_281, __A17_NET_279, __A17_NET_280, __A17_NET_280, __A17_NET_281, __A17_2__CCH10, GND, __A17_NET_281, __A17_2__RCH10_n, __A17_NET_277, CHWL14_n, __A17_2__WCH10_n, __A17_NET_304, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17058(__A17_NET_306, __A17_NET_304, __A17_NET_305, __A17_NET_305, __A17_NET_306, __A17_2__CCH10, GND, __A17_NET_306, __A17_2__RCH10_n, __A17_NET_301, CHWL16_n, __A17_2__WCH10_n, __A17_NET_303, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U17059(__A17_NET_306, RYWD14, __A17_NET_310, RYWD16, __A17_NET_294, __A17_2__WCH10_n, GND, __A17_2__CCH10, __A17_NET_295, WCH11_n, __A17_NET_300, CCH11, __A17_NET_298, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U17060(__A17_NET_310, __A17_NET_303, __A17_NET_309, __A17_NET_309, __A17_NET_310, __A17_2__CCH10, GND, __A17_NET_310, __A17_2__RCH10_n, __A17_NET_307, __A17_NET_296, GOJAM, __A17_NET_295, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U17061(__A17_NET_308, CHOR16_n_U17061_2,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17062(CH1213, __A17_NET_277, CH1214, __A17_NET_301, CH1414, __A17_NET_302, GND, __A17_NET_308, CH1316, __A17_NET_307, CH1416, __A17_NET_278, CH1413, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U17063(WCHG_n, XB0_n, CCHG_n, XT1_n, XB0_n, __A17_NET_296, GND, __A17_NET_297, CCHG_n, XT1_n, XB1_n, __A17_NET_294, XT1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U17064(__A17_NET_293, XT1_n, XB0_n, __A17_NET_298, __A17_NET_297, GOJAM, GND, XT1_n, XB1_n, __A17_NET_299,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U17065(__A17_NET_293, __A17_2__RCH10_n, __A17_NET_299, RCH11_n,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U18001(__A18_NET_189, MKEY1, __A18_NET_181, __A18_NET_181, __A18_NET_189, __A18_NET_182, GND, __A18_NET_189, __A18_1__RCH15_n, CH1501, MKEY2, __A18_NET_184, __A18_NET_194, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1) U18002(__A18_NET_189, __A18_NET_126, __A18_NET_194, __A18_NET_125, __A18_NET_192, __A18_NET_124, GND, __A18_NET_123, __A18_NET_193, __A18_NET_122, __A18_NET_121, __A18_NET_113, MAINRS, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U18003(__A18_NET_184, __A18_NET_194, __A18_NET_182, CH1502, __A18_NET_194, __A18_1__RCH15_n, GND, MKEY3, __A18_NET_179, __A18_NET_192, __A18_NET_192, __A18_NET_182, __A18_NET_179, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18004(CH1503, __A18_NET_192, __A18_1__RCH15_n, __A18_NET_193, MKEY4, __A18_NET_180, GND, __A18_NET_193, __A18_NET_182, __A18_NET_180, __A18_NET_193, __A18_1__RCH15_n, CH1504, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18005(__A18_NET_121, MKEY5, __A18_NET_120, __A18_NET_120, __A18_NET_121, __A18_NET_182, GND, __A18_NET_121, __A18_1__RCH15_n, CH1505, __A18_NET_123, __A18_NET_122, __A18_NET_188, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18006(__A18_NET_126, __A18_NET_125, __A18_NET_118, __A18_NET_116, __A18_1__F09D, __A18_NET_119, GND, KYRPT1, TPOR_n, __A18_NET_118, F09B_n, __A18_NET_187, __A18_NET_124, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U18007(__A18_NET_187, __A18_NET_116_U18007_2, __A18_NET_188, __A18_NET_116_U18007_4, __A18_NET_178, __A18_NET_99_U18007_6, GND, __A18_NET_99_U18007_8, __A18_NET_174, __A18_2__CNTOF9_U18007_10, __A18_NET_249, __A18_2__CNTOF9_U18007_12, __A18_NET_247, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U18008(__A18_NET_113, __A18_NET_182, __A18_NET_114, __A18_1__RCH15_n, __A18_NET_116, __A18_NET_127, GND, __A18_NET_105, NAVRST, __A18_NET_111, __A18_NET_105, __A18_1__RCH16_n, __A18_NET_112, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U18009(__A18_2__RRSYNC, __A18_NET_267, __A18_NET_257, __A18_NET_114, XT1_n, XB5_n, GND, __A18_NET_117, __A18_NET_119, __A18_NET_118, T05, T11, TPOR_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U18010(__A18_NET_117, __A18_1__F09A_n, __A18_NET_116, __A18_NET_182, __A18_NET_134,  , GND,  , __A18_1__F09A_n, __A18_NET_99, __A18_NET_111, __A18_NET_161, __A18_NET_100, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18011(__A18_NET_132, __A18_NET_127, __A18_NET_113, __A18_NET_134, __A18_NET_132, __A18_NET_133, GND, __A18_NET_134, KYRPT1, __A18_NET_133, XT1_n, XB6_n, __A18_NET_112, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U18012(__A18_NET_129, NKEY1, __A18_NET_128, __A18_NET_128, __A18_NET_129, __A18_NET_111, GND, __A18_NET_129, __A18_1__RCH16_n, CH1601, NKEY2, __A18_NET_130, __A18_NET_131, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U18013(__A18_NET_129, __A18_NET_110, __A18_NET_131, __A18_NET_109, __A18_NET_96, __A18_NET_108, GND, __A18_NET_107, __A18_NET_94, __A18_NET_106, __A18_NET_95, __A18_NET_162, __A18_NET_99, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U18014(__A18_NET_130, __A18_NET_131, __A18_NET_111, CH1602, __A18_NET_131, __A18_1__RCH16_n, GND, NKEY3, __A18_NET_97, __A18_NET_96, __A18_NET_96, __A18_NET_111, __A18_NET_97, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18015(CH1603, __A18_NET_96, __A18_1__RCH16_n, __A18_NET_94, NKEY4, __A18_NET_98, GND, __A18_NET_94, __A18_NET_111, __A18_NET_98, __A18_NET_94, __A18_1__RCH16_n, CH1604, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18016(__A18_NET_95, NKEY5, __A18_NET_93, __A18_NET_93, __A18_NET_95, __A18_NET_111, GND, __A18_NET_95, __A18_1__RCH16_n, CH1605, __A18_NET_107, __A18_NET_106, __A18_NET_174, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18017(__A18_NET_110, __A18_NET_109, __A18_NET_101, __A18_NET_99, __A18_1__F09D, __A18_NET_102, GND, KYRPT2, TPOR_n, __A18_NET_101, F09B_n, __A18_NET_178, __A18_NET_108, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U18018(__A18_NET_101, __A18_NET_100, __A18_NET_102, __A18_NET_103, __A18_NET_162, __A18_NET_105, GND, __A18_NET_103, __A18_NET_104, __A18_NET_161, __A18_NET_161, KYRPT2, __A18_NET_104, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18119(__A18_NET_164, WCH13_n, CHWL11_n, __A18_NET_165, __A18_NET_164, __A18_NET_163, GND, __A18_NET_165, CCH13, __A18_NET_163, __A18_NET_165, RCH13_n, CH1311, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0) U18120(SBYBUT, __A18_NET_158, F17A, __A18_1__F17A_n, F17B, __A18_1__F17B_n, GND, STNDBY_n, __A18_1__STNDBY, SBY, STNDBY_n, SBYLIT, __A18_NET_168, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18121(__A18_NET_155, __A18_1__F17A_n, __A18_NET_158, __A18_NET_157, __A18_NET_155, __A18_NET_156, GND, __A18_NET_157, __A18_NET_158, __A18_NET_156, __A18_1__F17B_n, __A18_NET_157, __A18_NET_159, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U18122(__A18_NET_170, __A18_NET_159, __A18_NET_160, __A18_NET_160, __A18_NET_170, __A18_NET_158, GND, __A18_NET_172, __A18_NET_167, __A18_NET_171, __A18_NET_171, __A18_NET_170, __A18_NET_167, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U18023( ,  , __A18_2__ACTV_n, RADRPT, CCH13, __A18_NET_263, GND, __A18_2__ADVCNT, F10A_n, __A18_NET_213, SB2_n,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18124(__A18_NET_166, __A18_NET_167, __A18_NET_170, __A18_NET_173, __A18_NET_167, __A18_1__STNDBY, GND, __A18_NET_173, __A18_NET_166, __A18_1__STNDBY, __A18_1__STNDBY, ALTEST, __A18_NET_168, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U18025(MRKRST, __A18_NET_135, __A18_NET_135, __A18_NET_146, __A18_NET_143, __A18_NET_151, GND, __A18_NET_149, __A18_NET_145, __A18_NET_150, __A18_NET_136, __A18_1__F08B_n, F08B, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U18026(__A18_NET_143, MARK, __A18_NET_169, __A18_NET_169, __A18_NET_143, __A18_NET_146, GND, MRKREJ, __A18_NET_144, __A18_NET_145, __A18_NET_145, __A18_NET_146, __A18_NET_144, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U18027(CH1606, __A18_NET_143, __A18_1__RCH16_n, CH1607, __A18_NET_145, __A18_1__RCH16_n, GND, __A18_NET_151, __A18_NET_149, __A18_NET_136, __A18_NET_137, __A18_NET_139, __A18_NET_138, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b0, 1'b1) U18028(__A18_NET_137, __A18_1__F09A_n, __A18_NET_136, __A18_NET_146, __A18_NET_142,  , GND,  , __A18_NET_231, RADRPT, __A18_2__ADVCNT, __A18_NET_251, __A18_NET_250, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18029(TPOR_n, __A18_NET_138, __A18_NET_138, __A18_NET_136, __A18_1__F09D, __A18_NET_139, GND, __A18_NET_260, __A18_NET_274, __A18_NET_273, __A18_NET_272, MKRPT, F09B_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18030(__A18_NET_140, __A18_NET_150, __A18_NET_135, __A18_NET_142, __A18_NET_140, __A18_NET_141, GND, __A18_NET_142, MKRPT, __A18_NET_141, __A18_NET_147, FS09_n, __A18_1__F09D, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1) U18031(__A18_1__F08B_n, __A18_NET_147, __A18_NET_220, __A18_NET_269, __A18_NET_208, __A18_NET_274, GND, __A18_NET_212, __A18_NET_207, __A18_NET_210, __A18_NET_206, __A18_NET_199, __A18_2__CNTOF9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U18032(__A18_NET_221, CHWL04_n, WCH13_n, __A18_2__ACTV_n, __A18_NET_221, __A18_NET_263, GND, RCH13_n, __A18_2__ACTV_n, CH1304, CHWL03_n, WCH13_n, __A18_NET_219, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18033(__A18_NET_220, __A18_NET_219, __A18_NET_208, __A18_NET_208, __A18_NET_220, CCH13, GND, RCH13_n, __A18_NET_220, CH1303, CHWL02_n, WCH13_n, __A18_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18034(__A18_NET_223, __A18_NET_222, __A18_NET_205, __A18_NET_205, __A18_NET_223, CCH13, GND, RCH13_n, __A18_NET_223, CH1302, CHWL01_n, WCH13_n, __A18_NET_217, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18035(__A18_NET_216, __A18_NET_217, __A18_NET_211, __A18_NET_211, __A18_NET_216, CCH13, GND, RCH13_n, __A18_NET_216, CH1301, F10A_n, SB0_n, __A18_2__F10AS0, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18036(__A18_NET_213, __A18_2__F10AS0, __A18_NET_214, __A18_NET_214, __A18_NET_213, __A18_2__ACTV_n, GND, __A18_NET_251, __A18_NET_253, __A18_NET_218, __A18_NET_250, __A18_NET_253, __A18_NET_228, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18037(__A18_NET_250, __A18_2__ADVCNT, __A18_NET_228, RADRPT, __A18_NET_250, __A18_NET_231, GND, __A18_NET_241, __A18_NET_254, __A18_NET_231, __A18_NET_230, __A18_NET_251, __A18_NET_218, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18038(__A18_NET_253, __A18_NET_228, __A18_NET_251, __A18_NET_229, __A18_NET_238, __A18_NET_254, GND, __A18_NET_241, __A18_NET_224, __A18_NET_230, __A18_NET_254, __A18_NET_224, __A18_NET_238, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b1) U18039(__A18_NET_254, __A18_NET_229, RADRPT, __A18_NET_231, __A18_NET_241,  , GND,  , __A18_NET_227, RADRPT, __A18_NET_229, __A18_NET_232, __A18_NET_234, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18040(__A18_NET_224, __A18_NET_238, __A18_NET_241, __A18_NET_227, __A18_NET_233, __A18_NET_234, GND, __A18_NET_232, __A18_NET_225, __A18_NET_226, __A18_NET_234, __A18_NET_225, __A18_NET_233, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18041(__A18_NET_234, __A18_NET_229, __A18_NET_235, __A18_NET_227, __A18_NET_198, __A18_NET_242, GND, __A18_NET_247, __A18_NET_224, __A18_NET_228, F10A, __A18_NET_232, __A18_NET_226, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U18042(__A18_NET_225, __A18_NET_233, __A18_NET_232, __A18_NET_196, __A18_NET_197, __A18_NET_235, GND, __A18_NET_242, __A18_NET_248, __A18_NET_198, __A18_NET_235, __A18_NET_248, __A18_NET_197, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U18043(__A18_NET_235, __A18_NET_196, RADRPT, __A18_NET_227, __A18_NET_242,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U18044(__A18_NET_248, __A18_NET_197, __A18_NET_242, __A18_NET_249, __A18_NET_197, __A18_NET_225, GND, __A18_2__ADVCNT, __A18_NET_195, __A18_NET_209, __A18_NET_205, __A18_NET_211, __A18_NET_265, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18045(__A18_NET_209, __A18_2__CNTOF9, __A18_NET_269, __A18_NET_209, F5BSB2_n, __A18_NET_207, GND, __A18_NET_206, F5BSB2_n, __A18_NET_209, __A18_NET_274, __A18_NET_195, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18046(__A18_NET_205, __A18_NET_216, __A18_NET_212, __A18_NET_211, __A18_NET_223, __A18_2__RRRARA, GND, __A18_2__LRXVEL, __A18_NET_211, __A18_NET_205, __A18_NET_210, __A18_2__RRRANG, __A18_NET_212, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18047(__A18_NET_210, __A18_NET_216, __A18_NET_210, __A18_NET_223, __A18_NET_211, __A18_2__LRZVEL, GND, __A18_2__LRRANG, __A18_NET_210, __A18_NET_223, __A18_NET_216, __A18_2__LRYVEL, __A18_NET_205, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U18048(__A18_NET_203, __A18_NET_199, GTSET_n, __A18_NET_202, __A18_NET_203, __A18_NET_204, GND, F5ASB2_n, __A18_NET_202, __A18_NET_256, __A18_NET_256, __A18_NET_200, __A18_NET_201, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18049(__A18_NET_202, RADRPT, __A18_NET_201, F09B, GOJAM, __A18_NET_200, GND, RADRPT, __A18_NET_270, __A18_NET_201, GTRST_n, __A18_NET_204, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0) U18050(TPOR_n, __A18_2__HERB, __A18_2__HERB, __A18_NET_270, __A18_NET_268, __A18_NET_267, GND, __A18_NET_266, RRIN1, __A18_NET_276, RRIN0, __A18_NET_275, LRIN1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U18051(__A18_NET_268, __A18_NET_265, __A18_NET_269, __A18_NET_259, __A18_NET_264, __A18_NET_262, GND, __A18_NET_261, __A18_NET_260, __A18_NET_258, __A18_NET_257, __A18_NET_274, __A18_2__LRSYNC, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U18052(__A18_NET_267, __A18_NET_266, __A18_NET_267, __A18_NET_276, __A18_NET_272, __A18_NET_261, GND, __A18_NET_262, __A18_NET_274, __A18_NET_275, __A18_NET_272, __A18_NET_264, __A18_NET_272, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U18053(LRIN0, __A18_NET_273, __A18_NET_263, __A18_NET_272, F09A, __A18_1__F09A_n, GND, RNRADP, __A18_NET_259, RNRADM, __A18_NET_258, __A18_NET_257, __A18_NET_256, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U18154(SBY, SBYREL_n,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U18155(__A18_NET_170, STOP,  ,  ,  ,  , GND,  ,  ,  ,  , __A18_NET_172, __A18_NET_165, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19001(__A19_NET_225, CA6_n, CXB0_n, __A19_NET_212, SHINC_n, T06_n, GND, __A19_NET_212, __A19_NET_213, __A19_1__SH3MS_n, __A19_1__SH3MS_n, CSG, __A19_NET_213, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1) U19002(__A19_NET_225, __A19_NET_214, __A19_NET_215, __A19_NET_209, __A19_NET_246, __A19_1__ALTSNC, GND, __A19_NET_235, __A19_NET_236, __A19_1__OTLNK0, __A19_NET_230, F5ASB0_n, __A19_1__F5ASB0, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19003(BR1, __A19_1__SH3MS_n, __A19_NET_214, __A19_1__SH3MS_n, BR1_n, __A19_NET_211, GND, __A19_NET_220, __A19_NET_221, CCH14, __A19_NET_226, __A19_NET_215, __A19_NET_214, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19004(__A19_NET_216, CHWL02_n, WCH14_n, __A19_NET_208, __A19_NET_216, __A19_NET_207, GND, __A19_NET_208, CCH14, __A19_NET_207, RCH14_n, __A19_NET_208, CH1402, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19005(__A19_1__ALT0, __A19_NET_209, __A19_NET_207, __A19_1__ALT1, __A19_NET_207, __A19_NET_210, GND, __A19_NET_209, __A19_NET_208, __A19_1__ALRT0, __A19_NET_208, __A19_NET_210, __A19_1__ALRT1, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19006(__A19_NET_210, __A19_NET_211, __A19_NET_218, __A19_NET_222, WCH14_n, CHWL03_n, GND, __A19_NET_222, __A19_NET_220, __A19_NET_221, __A19_NET_220, __A19_NET_226, __A19_NET_223, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19007(CH1403, RCH14_n, __A19_NET_223, __A19_NET_217, __A19_NET_224, __A19_NET_229, GND, __A19_NET_221, GTSET_n, __A19_NET_224, F5ASB2_n, __A19_NET_217, __A19_NET_218, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19008(__A19_NET_217, GOJAM, __A19_NET_219, GTSET, GOJAM, __A19_NET_226, GND, __A19_NET_246, __A19_NET_228, __A19_NET_226, __A19_NET_229, __A19_NET_229, GTONE, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U19009(__A19_NET_219, __A19_NET_218, __A19_NET_226, ALTM, F5ASB0_n, __A19_NET_219, GND, __A19_NET_226, __A19_NET_228, __A19_NET_227, __A19_NET_227, GTONE, __A19_NET_228, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U19010(__A19_NET_242, CHWL01_n, WCH14_n, __A19_NET_243, __A19_NET_242, __A19_NET_241, GND, GTSET_n, __A19_NET_243, __A19_NET_244, __A19_NET_244, __A19_NET_245, __A19_NET_248, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19011(__A19_NET_243, CCH14, __A19_NET_248, GTONE, GOJAM, __A19_NET_245, GND, __A19_NET_249, __A19_NET_247, GTSET, GOJAM, __A19_NET_241, __A19_NET_249, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19012(__A19_NET_232, F5ASB2_n, __A19_NET_248, __A19_NET_247, __A19_NET_232, __A19_NET_249, GND, F5ASB0_n, __A19_NET_247, OTLNKM, __A19_NET_241, __A19_NET_249, __A19_NET_231, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19013(CH1401, __A19_NET_231, RCH14_n, __A19_NET_230, __A19_NET_232, __A19_NET_234, GND, CA5_n, CXB7_n, __A19_NET_236, SB0_n, F05A_n, __A19_1__F5ASB0, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19014(BR1_n, __A19_1__SH3MS_n, __A19_NET_235, __A19_1__SH3MS_n, BR1, __A19_1__OTLNK1, GND, __A19_NET_176, __A19_NET_238, __A19_1__UPL0_n, __A19_1__BLKUPL, __A19_NET_234, __A19_NET_235, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19015(F5ASB2, F05A_n, SB2_n, __A19_1__F5BSB2, SB2_n, F05B_n, GND, __A19_1__XLNK0_n, __A19_NET_173, __A19_NET_169, __A19_1__XLNK1_n, __A19_NET_173, __A19_NET_172, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1) U19016(F5ASB2, F5ASB2_n, __A19_1__F5BSB2, F5BSB2_n, C45R, __A19_1__C45R_n, GND, __A19_NET_199, __A19_NET_198, __A19_NET_203, __A19_NET_202, __A19_1__UPL0_n, UPL0, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19017(__A19_1__BLKUPL, __A19_NET_238, __A19_NET_168, __A19_NET_165, __A19_NET_167, INLNKM, GND, INLNKP, __A19_NET_166, __A19_NET_165, __A19_NET_167, __A19_NET_177, __A19_1__UPL1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b0) U19018(__A19_NET_168, __A19_NET_176, __A19_NET_169, __A19_NET_166, __A19_NET_177, __A19_NET_172, GND, __A19_1__C45R_n, __A19_NET_182, __A19_NET_171, __A19_NET_171, __A19_NET_170, __A19_NET_182, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U19019(__A19_NET_178, __A19_NET_176, __A19_NET_177, __A19_NET_169, __A19_NET_172,  , GND,  , CA2_n, XB5_n, WOVR_n, OVF_n, T2P, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19020(__A19_NET_170, __A19_NET_171, __A19_NET_167, __A19_NET_167, __A19_NET_170, F04A, GND, BR1_n, __A19_1__C45R_n, UPRUPT, __A19_NET_170, __A19_NET_178, __A19_NET_180, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19021(__A19_NET_179, __A19_NET_180, __A19_NET_181, CH3311, __A19_NET_181, RCH33_n, GND, RCH33_n, __A19_1__BLKUPL, CH3310, CHWL05_n, WCH13_n, __A19_NET_159, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19022(__A19_NET_173, __A19_NET_159, __A19_NET_238, __A19_NET_238, __A19_NET_173, CCH13, GND, __A19_NET_173, CCH13, CH1305, WCH13_n, CHWL06_n, __A19_NET_163, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19023(__A19_NET_164, __A19_NET_163, __A19_NET_165, __A19_NET_165, __A19_NET_164, CCH13, GND, __A19_NET_164, CCH13, CH1306, CA5_n, XB5_n, __A19_NET_198, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19024(__A19_NET_179, CCH33, CCHG_n, XT3_n, XB3_n, CCH33, GND, __A19_NET_161, __A19_NET_196, __A19_NET_200, CCH14, __A19_NET_181, GOJAM, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19025(__A19_NET_194, __A19_NET_199, POUT_n, __A19_NET_197, __A19_NET_199, MOUT_n, GND, __A19_NET_199, ZOUT_n, __A19_NET_200, __A19_NET_162, __A19_NET_161, __A19_NET_196, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19026(__A19_NET_162, WCH14_n, CHWL04_n, CH1404, RCH14_n, __A19_NET_196, GND, __A19_NET_196, F5ASB2_n, THRSTD, __A19_NET_194, __A19_NET_195, __A19_NET_205, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19027(__A19_NET_195, __A19_NET_205, __A19_NET_196, __A19_NET_206, __A19_NET_197, __A19_NET_204, GND, __A19_NET_206, __A19_NET_196, __A19_NET_204, __A19_NET_205, F5ASB0_n, __A19_1__THRSTp, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19028(__A19_1__THRSTm, __A19_NET_206, F5ASB0_n, __A19_NET_202, CA5_n, XB6_n, GND, __A19_NET_203, POUT_n, __A19_NET_184, WCH14_n, CHWL05_n, __A19_NET_189, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19029(__A19_NET_186, __A19_NET_203, MOUT_n, __A19_NET_188, __A19_NET_203, ZOUT_n, GND, __A19_NET_189, __A19_NET_201, __A19_NET_190, RCH14_n, __A19_NET_190, CH1405, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19030(__A19_NET_190, __A19_NET_188, __A19_NET_328, __A19_NET_278, CCH14, __A19_NET_319, GND, __A19_NET_282, SB1_n, __A19_NET_271, __A19_NET_272, __A19_NET_201, CCH14, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U19031(EMSD, __A19_NET_190, F5ASB2_n, __A19_NET_192, __A19_NET_184, __A19_NET_185, GND, __A19_NET_192, __A19_NET_190, __A19_NET_185, __A19_NET_186, __A19_NET_187, __A19_NET_193, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19032(__A19_NET_187, __A19_NET_193, __A19_NET_190, __A19_1__EMSp, __A19_NET_192, F5ASB0_n, GND, __A19_NET_193, F5ASB0_n, __A19_1__EMSm, CHWL09_n, WCH11_n, __A19_NET_316, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0) U19033(BLKUPL_n, __A19_1__BLKUPL, UPL1, __A19_1__UPL1_n, XLNK0, __A19_1__XLNK0_n, GND, __A19_1__XLNK1_n, XLNK1, OUTCOM, __A19_2__FF1109_n, ERRST, __A19_NET_312, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19034(__A19_2__FF1109_n, __A19_NET_316, __A19_NET_317, __A19_NET_317, __A19_2__FF1109_n, CCH11, GND, RCH11_n, __A19_2__FF1109_n, CH1109, CHWL10_n, WCH11_n, __A19_NET_330, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19035(__A19_2__FF1110_n, __A19_NET_330, __A19_NET_318, __A19_NET_318, __A19_2__FF1110_n, CCH11, GND, CAURST, __A19_NET_330, __A19_NET_312, RCH11_n, __A19_2__FF1110_n, CH1110, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U19036(__A19_2__FF1110_n, __A19_2__OT1110, __A19_2__FF1111_n, __A19_2__OT1111, __A19_2__FF1112_n, __A19_2__OT1112, GND, __A19_NET_286, __A19_NET_282, __A19_NET_281, __A19_NET_283, __A19_NET_285, __A19_NET_284, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19037(__A19_NET_314, CHWL11_n, WCH11_n, __A19_2__FF1111_n, __A19_NET_314, __A19_NET_315, GND, __A19_2__FF1111_n, CCH11, __A19_NET_315, RCH11_n, __A19_2__FF1111_n, CH1111, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19038(__A19_NET_325, CHWL12_n, WCH11_n, __A19_2__FF1112_n, __A19_NET_325, __A19_NET_326, GND, __A19_2__FF1112_n, CCH11, __A19_NET_326, RCH11_n, __A19_2__FF1112_n, CH1112, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U19039(__A19_NET_329, CHWL10_n, WCH14_n, __A19_NET_328, __A19_NET_329, __A19_NET_319, GND, RCH14_n, __A19_NET_328, CH1410, CHWL09_n, WCH14_n, __A19_NET_320, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19040(__A19_NET_321, __A19_NET_320, __A19_NET_287, __A19_NET_287, __A19_NET_321, CCH14, GND, RCH14_n, __A19_NET_321, CH1409, CHWL08_n, WCH14_n, __A19_NET_322, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19041(__A19_NET_323, __A19_NET_322, __A19_NET_271, __A19_NET_271, __A19_NET_323, CCH14, GND, RCH14_n, __A19_NET_323, CH1408, CHWL07_n, WCH14_n, __A19_NET_311, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19042(__A19_NET_272, __A19_NET_311, __A19_NET_270, __A19_NET_270, __A19_NET_272, CCH14, GND, RCH14_n, __A19_NET_272, CH1407, CHWL06_n, WCH14_n, __A19_NET_273, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19043(__A19_NET_275, __A19_NET_273, __A19_NET_274, __A19_NET_274, __A19_NET_275, CCH14, GND, RCH14_n, __A19_NET_275, CH1406, __A19_NET_328, F5ASB2_n, GYROD, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19044(SB1_n, __A19_NET_270, SB1_n, __A19_NET_323, __A19_NET_272, __A19_NET_284, GND, __A19_NET_254, __A19_NET_255, __A19_NET_279, __A19_NET_280, __A19_NET_283, __A19_NET_323, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19045(__A19_2__GYENAB, SB1_n, __A19_NET_275, __A19_2__GYXP, __A19_NET_287, __A19_NET_286, GND, __A19_NET_286, __A19_NET_321, __A19_2__GYXM, __A19_NET_287, __A19_NET_281, __A19_2__GYYP, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19046(__A19_2__GYYM, __A19_NET_281, __A19_NET_321, __A19_2__GYZP, __A19_NET_287, __A19_NET_285, GND, __A19_NET_285, __A19_NET_321, __A19_2__GYZM, CA4_n, XB7_n, __A19_NET_276, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0) U19047(__A19_NET_276, __A19_NET_277, __A19_NET_252, __A19_2__O44, F06B, __A19_2__F06B_n, GND, __A19_2__F07D_n, __A19_NET_266, __A19_2__F07C_n, __A19_NET_267, __A19_2__F7CSB1_n, __A19_NET_268, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19048(__A19_NET_279, POUT_n, __A19_NET_277, __A19_NET_280, MOUT_n, __A19_NET_277, GND, ZOUT_n, __A19_NET_277, __A19_NET_278, __A19_NET_328, __A19_NET_254, __A19_NET_255, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19049(__A19_2__GYRRST, F5ASB2_n, __A19_NET_255, __A19_2__GYRSET, F5ASB2_n, __A19_NET_254, GND, CHWL08_n, WCH13_n, __A19_NET_256, __A19_NET_256, __A19_NET_252, __A19_NET_257, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U19050(__A19_NET_252, __A19_NET_257, CCH13, CH1308, RCH13_n, __A19_NET_257, GND, WCH13_n, CHWL09_n, __A19_NET_251, __A19_NET_251, __A19_NET_250, __A19_NET_253, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U19051(__A19_NET_262, __A19_NET_261, __A19_NET_300, CH1309, RCH13_n, __A19_NET_253, GND, __A19_NET_253, __A19_2__F07D_n, __A19_NET_269, FS07_n, __A19_2__F06B_n, __A19_NET_266, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U19052(__A19_NET_267, __A19_2__F06B_n, FS07A, __A19_NET_268, __A19_2__F07C_n, SB1_n, GND, __A19_NET_269, __A19_NET_259, __A19_NET_258, __A19_NET_258, F07B, __A19_NET_259, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19053(SB2_n, __A19_NET_258, __A19_NET_253, CCH13, __A19_2__RHCGO, __A19_NET_250, GND, __A19_NET_265, __A19_NET_260, __A19_2__F07C_n, SB0_n, __A19_2__RHCGO, __A19_2__F07C_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0) U19054(__A19_NET_259, __A19_NET_260, SB2, __A19_2__CNTRSB_n, F10B, __A19_2__F10B_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19055(SIGNX, __A19_2__F07C_n, SIGNY, __A19_2__F07C_n, __A19_2__F7CSB1_n, __A19_NET_263, GND, __A19_NET_264, SIGNZ, __A19_2__F07C_n, __A19_2__F7CSB1_n, __A19_NET_261, __A19_2__F7CSB1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U19056(__A19_NET_300, __A19_NET_262, __A19_NET_265, __A19_NET_302, __A19_NET_263, __A19_NET_303, GND, __A19_NET_302, __A19_NET_265, __A19_NET_303, __A19_NET_264, __A19_NET_309, __A19_NET_304, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19057(__A19_NET_309, __A19_NET_304, __A19_NET_265, __A19_NET_299, BMGXP, __A19_NET_310, GND, BMGXM, __A19_NET_301, __A19_NET_289, BMGYP, __A19_NET_305, __A19_NET_290, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19058(F5ASB2_n, __A19_NET_262, F5ASB2_n, __A19_NET_300, GATEX_n, __A19_NET_301, GND, __A19_NET_305, F5ASB2_n, __A19_NET_302, GATEY_n, __A19_NET_310, GATEX_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19059(F5ASB2_n, __A19_NET_303, F5ASB2_n, __A19_NET_304, GATEZ_n, __A19_NET_307, GND, __A19_NET_308, F5ASB2_n, __A19_NET_309, GATEZ_n, __A19_NET_306, GATEY_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19060(__A19_NET_291, BMGYM, __A19_NET_306, __A19_NET_292, BMGZP, __A19_NET_307, GND, BMGZM, __A19_NET_308, __A19_NET_293, __A19_2__O44, __A19_NET_299, BMAGXP, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19061(BMAGXM, __A19_2__O44, __A19_NET_289, BMAGYP, __A19_2__O44, __A19_NET_290, GND, __A19_2__O44, __A19_NET_291, BMAGYM, __A19_2__O44, __A19_NET_292, BMAGZP, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U19062(BMAGZM, __A19_2__O44, __A19_NET_293, T1P, __A19_2__CNTRSB_n, __A19_2__F10B_n, GND, __A19_2__F10B_n, __A19_2__CNTRSB_n, T3P, F10A_n, __A19_2__CNTRSB_n, T5P, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U19063(FS10, F09B_n, __A19_2__F06B_n, T6ON_n, __A19_2__CNTRSB_n, T6P, GND,  ,  ,  ,  , T4P, __A19_2__CNTRSB_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20001(__A20_NET_148, CDUXP, __A20_NET_145, __A20_NET_145, __A20_NET_148, __A20_1__C1R, GND, CDUXM, __A20_NET_146, __A20_NET_144, __A20_NET_144, __A20_1__C1R, __A20_NET_146, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U20002(BKTF_n, __A20_NET_175, RSSB, __A20_NET_173, __A20_NET_171, __CG11, GND, __CG21, __A20_NET_161, __A20_NET_132, RSSB, __A20_NET_121, BKTF_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20003(__A20_NET_143, __A20_NET_145, __A20_NET_146, __A20_NET_147, __A20_NET_175, __A20_NET_143, GND, __A20_NET_147, __A20_NET_142, __A20_NET_150, __A20_NET_150, __A20_1__C1R, __A20_NET_142, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20004(C32A, __CG22, __A20_NET_150, __A20_NET_139, CDUYP, __A20_NET_134, GND, __A20_NET_139, __A20_1__C2R, __A20_NET_134, CDUYM, __A20_NET_135, __A20_NET_140, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20005(__A20_NET_173, CA3_n, __A20_NET_148, CA3_n, CXB2_n, C32P, GND, C32M, __A20_NET_144, CA3_n, CXB2_n, __A20_1__C1R, CXB2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20006(__A20_NET_135, __A20_NET_140, __A20_1__C2R, __A20_NET_136, __A20_NET_134, __A20_NET_135, GND, __A20_NET_175, __A20_NET_136, __A20_NET_137, __A20_NET_137, __A20_NET_170, __A20_NET_138, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20007(__A20_NET_170, __A20_NET_138, __A20_1__C2R, __A20_NET_165, T2P, __A20_NET_172, GND, __A20_NET_165, __A20_1__C3R, __A20_NET_172, __A20_NET_175, __A20_NET_165, __A20_NET_167, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20008(__A20_NET_173, CA3_n, __A20_NET_139, CA3_n, CXB3_n, C33P, GND, C33M, __A20_NET_140, CA3_n, CXB3_n, __A20_1__C2R, CXB3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20009(__CG22, __A20_NET_142, __CG22, __A20_NET_142, __A20_NET_170, __A20_NET_171, GND, __A20_1__C3R, __A20_NET_173, CA2_n, CXB4_n, C33A, __A20_NET_138, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U20010(__A20_NET_166, __A20_NET_167, __A20_NET_168, __A20_NET_168, __A20_NET_166, __A20_1__C3R, GND, GND, __A20_NET_166, C24A, T1P, __A20_NET_177, __A20_NET_176, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20011(__A20_NET_177, __A20_NET_176, __A20_1__C4R, __A20_NET_156, __A20_NET_175, __A20_NET_176, GND, __A20_NET_156, __A20_NET_155, __A20_NET_157, __A20_NET_157, __A20_1__C4R, __A20_NET_155, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20012(__A20_NET_173, CA2_n, GND, __A20_NET_168, __A20_NET_157, C25A, GND, __A20_1__C5R, __A20_NET_173, CA2_n, CXB6_n, __A20_1__C4R, CXB5_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20013(__A20_NET_151, T3P, __A20_NET_158, __A20_NET_158, __A20_NET_151, __A20_1__C5R, GND, __A20_NET_175, __A20_NET_151, __A20_NET_152, __A20_NET_152, __A20_NET_160, __A20_NET_153, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20014(__A20_NET_160, __A20_NET_153, __A20_1__C5R, __A20_NET_103, CDUZP, __A20_NET_107, GND, __A20_NET_103, __A20_1__C6R, __A20_NET_107, CDUZM, __A20_NET_105, __A20_NET_104, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U20015(C26A, GND, __A20_NET_168, __A20_NET_155, __A20_NET_153,  , GND,  , GND, __A20_NET_168, __A20_NET_155, __A20_NET_160, __A20_NET_161, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20016(__A20_NET_105, __A20_NET_104, __A20_1__C6R, __A20_NET_100, __A20_NET_107, __A20_NET_105, GND, __A20_NET_121, __A20_NET_100, __A20_NET_101, __A20_NET_101, __A20_NET_98, __A20_NET_102, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20017(__A20_NET_98, __A20_NET_102, __A20_1__C6R, C34A, __CG11, __A20_NET_102, GND, TRNP, __A20_NET_97, __A20_NET_93, __A20_NET_93, __A20_1__C7R, __A20_NET_97, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20018(__A20_NET_132, CA3_n, __A20_NET_103, CA3_n, CXB4_n, C34P, GND, C34M, __A20_NET_104, CA3_n, CXB4_n, __A20_1__C6R, CXB4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20019(__A20_NET_92, TRNM, __A20_NET_94, __A20_NET_94, __A20_NET_92, __A20_1__C7R, GND, __A20_NET_97, __A20_NET_94, __A20_NET_96, __A20_NET_121, __A20_NET_96, __A20_NET_90, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20020(__A20_NET_91, __A20_NET_90, __A20_NET_99, __A20_NET_99, __A20_NET_91, __A20_1__C7R, GND, T4P, __A20_NET_125, __A20_NET_122, __A20_NET_122, __A20_1__C8R, __A20_NET_125, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20021(__A20_NET_132, CA3_n, __A20_NET_93, CA3_n, CXB5_n, C35P, GND, C35M, __A20_NET_92, CA3_n, CXB5_n, __A20_1__C7R, CXB5_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20022(__CG11, __A20_NET_98, __CG11, __A20_NET_98, __A20_NET_99, __A20_NET_115, GND, __A20_1__C8R, __A20_NET_132, CA2_n, CXB7_n, C35A, __A20_NET_91, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U20023(__A20_NET_115, __CG12, __A20_NET_120, __CG22, __A20_NET_203, __CG14, GND, __CG24, __A20_NET_208,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20024(__A20_NET_124, __A20_NET_121, __A20_NET_122, __A20_NET_123, __A20_NET_124, __A20_NET_113, GND, __A20_NET_123, __A20_1__C8R, __A20_NET_113, __CG21, __A20_NET_123, C27A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20025(__A20_NET_127, T5P, __A20_NET_131, __A20_NET_131, __A20_NET_127, __A20_1__C9R, GND, __A20_NET_121, __A20_NET_127, __A20_NET_128, __A20_NET_128, __A20_NET_129, __A20_NET_130, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20026(__A20_NET_129, __A20_NET_130, __A20_1__C9R, __A20_NET_108, T6P, __A20_NET_112, GND, __A20_NET_108, __A20_1__C10R, __A20_NET_112, __A20_NET_121, __A20_NET_108, __A20_NET_110, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20027(__A20_NET_132, CA3_n, __CG21, __A20_NET_113, __A20_NET_130, C30A, GND, __A20_1__C10R, __A20_NET_132, CA3_n, CXB1_n, __A20_1__C9R, CXB0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20028(__A20_NET_109, __A20_NET_110, __A20_NET_111, __A20_NET_111, __A20_NET_109, __A20_1__C10R, GND, __A20_NET_198, __A20_NET_196, __A20_NET_199, __A20_NET_199, __A20_2__C10R, __A20_NET_196, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U20029(C31A, __CG21, __A20_NET_113, __A20_NET_129, __A20_NET_109,  , GND,  , __CG21, __A20_NET_113, __A20_NET_129, __A20_NET_111, __A20_NET_120, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20030(__A20_NET_235, PIPYP, __A20_NET_231, __A20_NET_231, __A20_NET_235, __A20_2__C1R, GND, PIPYM, __A20_NET_232, __A20_NET_236, __A20_NET_236, __A20_2__C1R, __A20_NET_232, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U20031(BKTF_n, __A20_NET_263, RSSB, __A20_NET_261, __A20_NET_259, CG13, GND, CG23, __A20_NET_251, __A20_NET_220, RSSB, __A20_NET_209, BKTF_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20032(__A20_NET_233, __A20_NET_231, __A20_NET_232, __A20_NET_234, __A20_NET_263, __A20_NET_233, GND, __A20_NET_234, __A20_NET_230, __A20_NET_237, __A20_NET_237, __A20_2__C1R, __A20_NET_230, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20033(C40A, __CG14, __A20_NET_237, __A20_NET_227, PIPZP, __A20_NET_223, GND, __A20_NET_227, __A20_2__C2R, __A20_NET_223, PIPZM, __A20_NET_224, __A20_NET_228, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20034(__A20_NET_261, CA4_n, __A20_NET_235, CA4_n, CXB0_n, C40P, GND, C40M, __A20_NET_236, CA4_n, CXB0_n, __A20_2__C1R, CXB0_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20035(__A20_NET_224, __A20_NET_228, __A20_2__C2R, __A20_NET_225, __A20_NET_223, __A20_NET_224, GND, __A20_NET_263, __A20_NET_225, __A20_NET_226, __A20_NET_226, __A20_NET_258, __A20_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20036(__A20_NET_258, __A20_NET_222, __A20_2__C2R, __A20_NET_254, TRUND, __A20_NET_260, GND, __A20_NET_254, __A20_2__C3R, __A20_NET_260, __A20_NET_263, __A20_NET_254, __A20_NET_256, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20037(__A20_NET_261, CA4_n, __A20_NET_227, CA4_n, CXB1_n, C41P, GND, C41M, __A20_NET_228, CA4_n, CXB1_n, __A20_2__C2R, CXB1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20038(__CG14, __A20_NET_230, __CG14, __A20_NET_230, __A20_NET_258, __A20_NET_259, GND, __A20_2__C3R, __A20_NET_261, CA5_n, CXB3_n, C41A, __A20_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U20039(__A20_NET_255, __A20_NET_256, __A20_NET_246, __A20_NET_246, __A20_NET_255, __A20_2__C3R, GND, __CG24, __A20_NET_255, C53A, SHAFTD, __A20_NET_265, __A20_NET_264, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20040(__A20_NET_265, __A20_NET_264, __A20_2__C4R, __A20_NET_245, __A20_NET_263, __A20_NET_264, GND, __A20_NET_245, __A20_NET_244, __A20_NET_243, __A20_NET_243, __A20_2__C4R, __A20_NET_244, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20041(__A20_NET_261, CA5_n, __CG24, __A20_NET_246, __A20_NET_243, C54A, GND, __A20_2__C5R, __A20_NET_261, CA5_n, CXB5_n, __A20_2__C4R, CXB4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20042(__A20_NET_239, THRSTD, __A20_NET_247, __A20_NET_247, __A20_NET_239, __A20_2__C5R, GND, __A20_NET_263, __A20_NET_239, __A20_NET_240, __A20_NET_240, __A20_NET_250, __A20_NET_241, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20043(__A20_NET_250, __A20_NET_241, __A20_2__C5R, __A20_NET_195, SHAFTP, __A20_NET_194, GND, __A20_NET_195, __A20_2__C6R, __A20_NET_194, SHAFTM, __A20_NET_191, __A20_NET_192, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U20044(C55A, __CG24, __A20_NET_246, __A20_NET_244, __A20_NET_241,  , GND,  , __CG24, __A20_NET_246, __A20_NET_244, __A20_NET_250, __A20_NET_251, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20045(__A20_NET_191, __A20_NET_192, __A20_2__C6R, __A20_NET_188, __A20_NET_194, __A20_NET_191, GND, __A20_NET_209, __A20_NET_188, __A20_NET_189, __A20_NET_189, __A20_NET_186, __A20_NET_190, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U20046(__A20_NET_186, __A20_NET_190, __A20_2__C6R, C36A, __CG12, __A20_NET_190, GND, PIPXP, __A20_NET_185, __A20_NET_181, __A20_NET_181, __A20_2__C7R, __A20_NET_185, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20047(__A20_NET_220, CA3_n, __A20_NET_195, CA3_n, CXB6_n, C36P, GND, C36M, __A20_NET_192, CA3_n, CXB6_n, __A20_2__C6R, CXB6_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20048(__A20_NET_180, PIPXM, __A20_NET_182, __A20_NET_182, __A20_NET_180, __A20_2__C7R, GND, __A20_NET_185, __A20_NET_182, __A20_NET_184, __A20_NET_209, __A20_NET_184, __A20_NET_178, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U20049(__A20_NET_179, __A20_NET_178, __A20_NET_187, __A20_NET_187, __A20_NET_179, __A20_2__C7R, GND, CDUXD, __A20_NET_213, __A20_NET_210, __A20_NET_210, __A20_2__C8R, __A20_NET_213, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20050(__A20_NET_220, CA3_n, __A20_NET_181, CA3_n, CXB7_n, C37P, GND, C37M, __A20_NET_180, CA3_n, CXB7_n, __A20_2__C7R, CXB7_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20051(__CG12, __A20_NET_186, __CG12, __A20_NET_186, __A20_NET_187, __A20_NET_203, GND, __A20_2__C8R, __A20_NET_220, CA5_n, CXB0_n, C37A, __A20_NET_179, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U20052(__A20_NET_212, __A20_NET_209, __A20_NET_210, __A20_NET_211, __A20_NET_212, __A20_NET_201, GND, __A20_NET_211, __A20_2__C8R, __A20_NET_201, CG26, __A20_NET_211, C50A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U20053(__A20_NET_215, CDUYD, __A20_NET_219, __A20_NET_219, __A20_NET_215, __A20_2__C9R, GND, __A20_NET_209, __A20_NET_215, __A20_NET_216, __A20_NET_216, __A20_NET_217, __A20_NET_218, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U20054(__A20_NET_217, __A20_NET_218, __A20_2__C9R, __A20_NET_197, CDUZD, __A20_NET_200, GND, __A20_NET_197, __A20_2__C10R, __A20_NET_200, __A20_NET_209, __A20_NET_197, __A20_NET_198, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U20055(__A20_NET_220, CA5_n, CG26, __A20_NET_201, __A20_NET_218, C51A, GND, __A20_2__C10R, __A20_NET_220, CA5_n, CXB2_n, __A20_2__C9R, CXB1_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U20056(C52A, CG26, __A20_NET_201, __A20_NET_217, __A20_NET_199,  , GND,  , CG26, __A20_NET_201, __A20_NET_217, __A20_NET_196, __A20_NET_208, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21001(__A21_NET_205, C25A, C27A, C31A, C33A,  , GND,  , C35A, C37A, C41A, __A21_1__C43A, __A21_NET_204, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21002(__A21_NET_205, __A21_NET_152_U21002_2, __A21_NET_204, __A21_NET_152_U21002_4, __A21_NET_199, __A21_NET_152_U21002_6, GND, __A21_NET_152_U21002_8, __A21_NET_200, __A21_NET_153_U21002_10, __A21_NET_203, __A21_NET_153_U21002_12, __A21_NET_219, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21003(__A21_NET_199, __A21_1__C45A, __A21_1__C47A, C51A, C53A,  , GND,  , C26A, C27A, C32A, C33A, __A21_NET_203, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U21004(__A21_NET_200, C55A, __A21_1__C57A, __A21_NET_225, __A21_1__C56A, __A21_1__C57A, GND, __A21_1__30SUM, __A21_1__C60A, __A21_NET_188, __A21_1__50SUM, __A21_1__C60A, __A21_NET_185, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21005(__A21_NET_219, C36A, C37A, __A21_1__C42A, __A21_1__C43A,  , GND,  , __A21_1__C46A, __A21_1__C47A, C52A, C53A, __A21_NET_224, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21006(__A21_NET_224, __A21_NET_153_U21006_2, __A21_NET_225, __A21_NET_153_U21006_4, __A21_NET_212, __A21_NET_147_U21006_6, GND, __A21_NET_147_U21006_8, __A21_NET_215, __A21_NET_147_U21006_10, __A21_NET_216, __A21_NET_147_U21006_12, __A21_NET_178, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21007(__A21_NET_212, C24A, C25A, C26A, C27A,  , GND,  , C34A, C35A, C36A, C37A, __A21_NET_215, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21008(__A21_NET_216, __A21_1__C44A, __A21_1__C45A, __A21_1__C46A, __A21_1__C47A,  , GND,  , C54A, C55A, __A21_1__C56A, __A21_1__C57A, __A21_NET_178, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21009(__A21_NET_179, C30A, C31A, C32A, C33A,  , GND,  , C34A, C35A, C36A, C37A, __A21_NET_184, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21010(__A21_NET_179, __A21_1__32004K_U21010_2, __A21_NET_184, __A21_1__32004K_U21010_4, __A21_NET_168, __A21_NET_173_U21010_6, GND, __A21_NET_173_U21010_8, __A21_NET_172, __A21_NET_146_U21010_10, __A21_NET_174, __A21_NET_146_U21010_12, __A21_NET_188, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U21011(__A21_1__32004K, __A21_1__30SUM, __A21_NET_173, __A21_1__50SUM, DINC, DINC_n, GND, CXB0_n, XB0, CXB1_n, XB1, CXB2_n, XB2, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21012(__A21_NET_168, C50A, C51A, C52A, C53A,  , GND,  , C54A, C55A, __A21_1__C56A, __A21_1__C57A, __A21_NET_172, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21013(__A21_NET_174, C24A, C25A, C26A, C27A,  , GND,  , C40A, C41A, __A21_1__C42A, __A21_1__C43A, __A21_NET_193, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21014(__A21_NET_193, __A21_NET_187_U21014_2, __A21_NET_194, __A21_NET_187_U21014_4, __A21_NET_185, __A21_NET_187_U21014_6, GND, __A21_NET_229_U21014_8, __A21_NET_228, __A21_NET_229_U21014_10, __A21_NET_227, __A21_NET_229_U21014_12, __A21_NET_226, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21015(__A21_NET_194, __A21_1__C44A, __A21_1__C45A, __A21_1__C46A, __A21_1__C47A,  , GND,  , __A21_1__C45M, __A21_1__C46M, __A21_1__C57A, __A21_1__C60A, __A21_NET_148, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U21016(__A21_NET_151, __A21_1__30SUM, __A21_1__50SUM, CAD1, __A21_1__RSCT_n, __A21_NET_152, GND, __A21_1__RSCT_n, __A21_NET_153, CAD2, __A21_1__RSCT_n, __A21_NET_147, CAD3, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U21017(CAD4, __A21_1__RSCT_n, __A21_NET_151, CAD5, __A21_1__RSCT_n, __A21_NET_146, GND, __A21_1__RSCT_n, __A21_NET_187, CAD6, __A21_1__C45P, __A21_1__C46P, __A21_NET_149, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21018(C31A, __A21_1__C47A, C51A, C52A, C53A, __A21_NET_227, GND, __A21_NET_226, C54A, C55A, __A21_1__C56A, __A21_NET_228, C50A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U21019(__A21_NET_156, INCSET_n, __A21_NET_148, __A21_NET_157, INCSET_n, __A21_NET_149, GND, INCSET_n, __A21_NET_229, __A21_NET_154, __A21_NET_156, __A21_1__SHINC, SHINC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21020(__A21_1__SHINC, SHINC_n, T12A, SHANC_n, __A21_NET_157, __A21_1__SHANC, GND, SHANC_n, T12A, __A21_1__SHANC, __A21_NET_154, DINC, __A21_1__DINCNC_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21021(DINC, __A21_1__DINCNC_n, T12A, __A21_NET_133, INCSET_n, __A21_NET_141, GND, __A21_NET_133, PINC, __A21_1__PINC_n, __A21_1__PINC_n, T12, PINC, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21022(__A21_NET_136, C24A, C25A, C26A, C27A,  , GND,  , C30A, C37P, C40P, C41P, __A21_NET_140, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21023(__A21_NET_136, __A21_NET_141_U21023_2, __A21_NET_140, __A21_NET_141_U21023_4, __A21_NET_134, __A21_NET_141_U21023_6, GND, __A21_NET_145_U21023_8, __A21_NET_144, __A21_NET_145_U21023_10, __A21_NET_142, __A21_NET_159_U21023_12, __A21_NET_164, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21024(__A21_1__C42P, __A21_1__C43P, __A21_1__C42M, __A21_1__C43M, __A21_1__C44M, __A21_NET_144, GND, __A21_NET_142, C37M, C40M, C41M, __A21_NET_134, __A21_1__C44P, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21025(__A21_NET_143, INCSET_n, __A21_NET_145, __A21_1__MINC_n, __A21_NET_143, MINC, GND, __A21_1__MINC_n, T12A, MINC, C35P, C36P, __A21_NET_160, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21026(C32P, C33P, C32M, C33M, C34M, __A21_NET_161, GND,  ,  ,  ,  , __A21_NET_164, C34P, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U21027(__A21_NET_160, __A21_NET_159_U21027_2, __A21_NET_161, __A21_NET_162_U21027_4, __A21_NET_163, __A21_NET_162_U21027_6, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21028(__A21_NET_166, INCSET_n, __A21_NET_159, __A21_1__PCDU_n, __A21_NET_166, PCDU, GND, __A21_1__PCDU_n, T12A, PCDU, C35M, C36M, __A21_NET_163, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21029(__A21_NET_165, INCSET_n, __A21_NET_162, __A21_1__MCDU_n, __A21_NET_165, MCDU, GND, __A21_1__MCDU_n, T12A, MCDU, __A21_NET_249, __A21_3__C43R, __A21_NET_252, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21030(__A21_NET_300, BMAGXP, __A21_NET_305, __A21_NET_305, __A21_NET_300, __A21_3__C42R, GND, BMAGXM, __A21_NET_304, __A21_NET_302, __A21_NET_302, __A21_3__C42R, __A21_NET_304, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0) U21031(BKTF_n, __A21_NET_301, RSSB, __A21_NET_276, __A21_NET_262, __A21_3__CG15, GND, CTROR, CTROR_n, __A21_NET_244, RSSB, __A21_NET_241, BKTF_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21032(__A21_NET_306, __A21_NET_305, __A21_NET_304, __A21_NET_307, __A21_NET_301, __A21_NET_306, GND, __A21_NET_307, __A21_NET_261, __A21_NET_308, __A21_NET_308, __A21_3__C42R, __A21_NET_261, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21033(__A21_1__C42A, CG13, __A21_NET_308, __A21_NET_249, BMAGYP, __A21_NET_252, GND, __A21_1__SHINC, __A21_1__SHANC, SHIFT_n, BMAGYM, __A21_NET_253, __A21_NET_250, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21034(__A21_NET_276, CA4_n, __A21_NET_300, CA4_n, CXB2_n, __A21_1__C42P, GND, __A21_1__C42M, __A21_NET_302, CA4_n, CXB2_n, __A21_3__C42R, CXB2_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21035(__A21_NET_253, __A21_NET_250, __A21_3__C43R, __A21_NET_254, __A21_NET_252, __A21_NET_253, GND, __A21_NET_301, __A21_NET_254, __A21_NET_256, __A21_NET_256, __A21_NET_255, __A21_NET_251, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21036(__A21_NET_255, __A21_NET_251, __A21_3__C43R, __A21_NET_264, EMSD, __A21_NET_263, GND, __A21_NET_264, __A21_3__C56R, __A21_NET_263, __A21_NET_301, __A21_NET_264, __A21_NET_258, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21037(__A21_NET_276, CA4_n, __A21_NET_249, CA4_n, CXB3_n, __A21_1__C43P, GND, __A21_1__C43M, __A21_NET_250, CA4_n, CXB3_n, __A21_3__C43R, CXB3_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21038(CG13, __A21_NET_261, CG13, __A21_NET_261, __A21_NET_255, __A21_NET_262, GND, __A21_3__C56R, __A21_NET_276, CA5_n, CXB6_n, __A21_1__C43A, __A21_NET_251, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U21039(__A21_NET_257, __A21_NET_258, __A21_NET_236, __A21_NET_236, __A21_NET_257, __A21_3__C56R, GND, CG23, __A21_NET_257, __A21_1__C56A, OTLNKM, __A21_NET_259, __A21_NET_260, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21040(__A21_NET_259, __A21_NET_260, __A21_3__C57R, __A21_NET_238, __A21_NET_301, __A21_NET_260, GND, __A21_NET_238, __A21_NET_245, __A21_NET_237, __A21_NET_237, __A21_3__C57R, __A21_NET_245, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21041(__A21_NET_276, CA5_n, CG23, __A21_NET_236, __A21_NET_237, __A21_1__C57A, GND, __A21_3__C60R, __A21_NET_276, CA6_n, CXB0_n, __A21_3__C57R, CXB7_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U21042(__A21_NET_234, ALTM, __A21_NET_239, __A21_NET_239, __A21_NET_234, __A21_3__C60R, GND, __A21_NET_301, __A21_NET_234, __A21_NET_235, __A21_NET_235, __A21_NET_233, __A21_NET_232, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21043(__A21_NET_233, __A21_NET_232, __A21_3__C60R, __A21_NET_288, BMAGZP, __A21_NET_246, GND, __A21_NET_288, __A21_3__C44R, __A21_NET_246, BMAGZM, __A21_NET_247, __A21_NET_248, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U21044(__A21_1__C60A, CG23, __A21_NET_236, __A21_NET_245, __A21_NET_232,  , GND,  , CG23, __A21_NET_236, __A21_NET_245, __A21_NET_233, CTROR_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21045(__A21_NET_247, __A21_NET_248, __A21_3__C44R, __A21_NET_240, __A21_NET_246, __A21_NET_247, __A21_NET_71, __A21_NET_241, __A21_NET_240, __A21_NET_243, __A21_NET_243, __A21_NET_292, __A21_NET_242, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U21046(__A21_NET_292, __A21_NET_242, __A21_3__C44R, __A21_1__C44A, __A21_3__CG15, __A21_NET_242, GND, INLNKP, __A21_NET_283, __A21_NET_289, __A21_NET_289, C45R, __A21_NET_283, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21047(__A21_NET_244, CA4_n, __A21_NET_288, CA4_n, CXB4_n, __A21_1__C44P, GND, __A21_1__C44M, __A21_NET_248, CA4_n, CXB4_n, __A21_3__C44R, CXB4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21048(__A21_NET_282, INLNKM, __A21_NET_281, __A21_NET_281, __A21_NET_282, C45R, GND, __A21_NET_283, __A21_NET_281, __A21_NET_284, __A21_NET_241, __A21_NET_284, __A21_NET_287, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U21049(__A21_NET_286, __A21_NET_287, __A21_NET_285, __A21_NET_285, __A21_NET_286, C45R, GND, RNRADP, __A21_NET_290, __A21_NET_275, __A21_NET_275, __A21_3__C46R, __A21_NET_290, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21050(__A21_NET_244, CA4_n, __A21_NET_289, CA4_n, CXB5_n, __A21_1__C45P, GND, __A21_1__C45M, __A21_NET_282, CA4_n, CXB5_n, C45R, CXB5_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21051(__A21_3__CG15, __A21_NET_292, __A21_3__CG15, __A21_NET_292, __A21_NET_285, __A21_NET_277, GND, __A21_3__C46R, __A21_NET_244, CA4_n, CXB6_n, __A21_1__C45A, __A21_NET_286, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U21052(__A21_NET_277, __A21_3__CG16, __A21_NET_278, CG26, XB3, CXB3_n, GND, CXB4_n, XB4, CXB5_n, XB5, CXB6_n, XB6, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b1) U21053(__A21_NET_273, __A21_NET_241, __A21_NET_280, __A21_NET_272, __A21_NET_273, __A21_NET_271, GND, __A21_NET_272, __A21_3__C46R, __A21_NET_271, __A21_3__CG16, __A21_NET_272, __A21_1__C46A, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U21054(__A21_NET_274, RNRADM, __A21_NET_279, __A21_NET_279, __A21_NET_274, __A21_3__C46R, GND, __A21_NET_290, __A21_NET_279, __A21_NET_280, __A21_NET_269, __A21_NET_265, __A21_NET_268, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U21055(__A21_NET_265, __A21_NET_268, __A21_3__C47R, __A21_NET_267, GYROD, __A21_NET_266, GND, __A21_NET_267, __A21_3__C47R, __A21_NET_266, __A21_NET_241, __A21_NET_267, __A21_NET_269, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21056(__A21_NET_275, CA4_n, CA4_n, CXB6_n, __A21_NET_274, __A21_1__C46M, GND, __A21_3__C47R, __A21_NET_244, CA4_n, CXB7_n, __A21_1__C46P, CXB6_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U21057(__A21_3__CG16, __A21_NET_271, __A21_3__CG16, __A21_NET_271, __A21_NET_265, __A21_NET_278, GND,  ,  ,  ,  , __A21_1__C47A, __A21_NET_268, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U21058(XB7, CXB7_n, OCTAD2, CA2_n, OCTAD3, CA3_n, GND, CA4_n, OCTAD4, CA5_n, OCTAD5, CA6_n, OCTAD6, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U21059(SHIFT_n, SHIFT, RSCT, __A21_1__RSCT_n,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U22001(__A22_NET_128, __A22_1__DLKRPT, __A22_NET_127, DLKPLS, T10_n, __A22_NET_128, GND, __A22_NET_133, __A22_NET_124, __A22_1__DLKRPT, __A22_1__DLKRPT, __A22_NET_123, __A22_NET_124, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22002(__A22_NET_128, DRPRST, __A22_NET_133, __A22_1__DLKRPT, __A22_NET_123, __A22_NET_129, GND, __A22_1__ADVCTR, __A22_1__RDOUT_n, __A22_1__WDORDR, __A22_1__BSYNC_n, __A22_NET_127, GOJAM, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0) U22003(DKEND, __A22_NET_133, __A22_NET_133, __A22_1__END, DKSTRT, __A22_NET_132, GND, __A22_1__DLKCLR, __A22_NET_132, __A22_NET_111, __A22_NET_109, __A22_1__DKCTR1_n, __A22_NET_117, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U22004(__A22_NET_123, __A22_1__DLKRPT, __A22_NET_125, __A22_NET_125, __A22_NET_123, F10A, GND, __A22_NET_129, __A22_NET_131, __A22_NET_130, __A22_NET_130, CCH33, __A22_NET_131, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U22005(CH3312, RCH33_n, __A22_NET_131, __A22_NET_109, __A22_1__DLKCLR, __A22_1__ADVCTR, GND, __A22_1__DLKCLR, __A22_NET_112, __A22_1__RDOUT_n, __A22_1__RDOUT_n, __A22_1__END, __A22_NET_112, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U22006(__A22_1__1CNT, __A22_NET_111, __A22_NET_121, __A22_NET_111, __A22_NET_118, __A22_NET_122, GND, __A22_NET_116, __A22_NET_117, __A22_1__DLKCLR, __A22_NET_122, __A22_NET_121, __A22_NET_122, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b1) U22007(__A22_1__1CNT, __A22_NET_117, __A22_NET_121, __A22_NET_118, __A22_NET_122, __A22_NET_116, GND, __A22_NET_121, __A22_NET_116, __A22_NET_117, __A22_NET_146, __A22_NET_119, __A22_NET_120, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U22008(__A22_NET_116, __A22_1__DKCTR1, __A22_NET_146, __A22_1__DKCTR2_n, __A22_NET_147, __A22_1__DKCTR2, GND, __A22_1__DKCTR3_n, __A22_NET_137, __A22_1__DKCTR3, __A22_NET_138, __A22_1__DKCTR4_n, __A22_NET_144, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U22009(__A22_NET_120, __A22_NET_118, __A22_NET_119, __A22_NET_118, __A22_NET_150, __A22_NET_148, GND, __A22_NET_147, __A22_NET_146, __A22_1__DLKCLR, __A22_NET_148, __A22_NET_119, __A22_NET_148, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U22010(__A22_NET_150, __A22_NET_148, __A22_NET_147, __A22_NET_146, __A22_NET_119, __A22_NET_147, GND, __A22_NET_137, __A22_NET_151, __A22_NET_149, __A22_NET_152, __A22_NET_138, __A22_NET_139, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U22011(__A22_NET_149, __A22_NET_150, __A22_NET_151, __A22_NET_150, __A22_NET_139, __A22_NET_152, GND, __A22_NET_138, __A22_NET_137, __A22_1__DLKCLR, __A22_NET_152, __A22_NET_151, __A22_NET_152, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b1, 1'b0, 1'b1) U22012(__A22_NET_137, __A22_NET_151, __A22_NET_138, __A22_NET_135, __A22_NET_144, __A22_NET_136, GND, __A22_NET_143, __A22_NET_145, __A22_NET_140, __A22_NET_136, __A22_NET_145, __A22_NET_144, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U22013(__A22_NET_135, __A22_NET_139, __A22_NET_136, __A22_NET_139, __A22_NET_140, __A22_NET_143, GND, __A22_NET_145, __A22_NET_144, __A22_1__DLKCLR, __A22_NET_143, __A22_NET_136, __A22_NET_143, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1) U22014(__A22_NET_145, __A22_1__DKCTR4, __A22_NET_74, __A22_1__DKCTR5_n, __A22_NET_75, __A22_1__DKCTR5, GND, __A22_NET_85, __A22_1__BSYNC_n, __A22_NET_84, __A22_NET_83, __A22_NET_79, __A22_NET_84, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U22015(__A22_1__16CNT, __A22_NET_74, __A22_NET_141, __A22_1__32CNT, __A22_NET_142, __A22_NET_75, GND, __A22_NET_141, __A22_NET_75, __A22_NET_74, __A22_NET_85, __A22_NET_79, __A22_NET_82, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U22016(__A22_1__16CNT, __A22_NET_140, __A22_NET_141, __A22_NET_140, __A22_1__32CNT, __A22_NET_142, GND, __A22_NET_75, __A22_NET_74, __A22_1__DLKCLR, __A22_NET_142, __A22_NET_141, __A22_NET_142, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22017(__A22_NET_78, __A22_NET_82, __A22_NET_83, __A22_NET_83, __A22_NET_85, __A22_NET_78, GND, CHWL07_n, WCH13_n, __A22_NET_80, __A22_NET_81, __A22_NET_80, __A22_NET_64, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U22018(__A22_NET_81, CCH13, __A22_NET_64, CH1307, RCH13_n, __A22_NET_64, GND, __A22_1__DLKCLR, __A22_1__WDORDR, __A22_NET_60, __A22_NET_60, __A22_NET_82, __A22_1__WDORDR, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U22019(__A22_1__ORDRBT, __A22_NET_64, __A22_NET_60, __A22_NET_58, __A22_1__DKCTR5, __A22_1__DKCTR4, GND, __A22_1__DKCTR5, __A22_1__DKCTR4_n, __A22_NET_61, __A22_1__DKCTR4, __A22_1__DKCTR5_n, __A22_NET_69, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U22020(__A22_NET_58, __A22_1__HIGH0_n, __A22_NET_61, __A22_1__HIGH1_n, __A22_NET_69, __A22_1__HIGH2_n, GND, __A22_1__HIGH3_n, __A22_NET_71, __A22_1__LOW0_n, __A22_NET_67, __A22_1__LOW1_n, __A22_NET_66, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22021(__A22_NET_71, __A22_1__DKCTR4_n, __A22_1__DKCTR5_n, __A22_NET_103, CHWL16_n, WCH34_n, GND, __A22_NET_103, __A22_NET_104, __A22_NET_91, __A22_NET_91, CCH34, __A22_NET_104, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22022(__A22_1__DKCTR1, __A22_1__DKCTR2, __A22_1__DKCTR1_n, __A22_1__DKCTR2, __A22_1__DKCTR3, __A22_NET_66, GND, __A22_NET_68, __A22_1__DKCTR1, __A22_1__DKCTR2_n, __A22_1__DKCTR3, __A22_NET_67, __A22_1__DKCTR3, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U22023(__A22_NET_68, __A22_1__LOW2_n, __A22_NET_102, __A22_1__LOW3_n, __A22_NET_96, __A22_1__LOW4_n, GND, __A22_1__LOW5_n, __A22_NET_100, __A22_1__LOW6_n, __A22_NET_107, __A22_1__LOW7_n, __A22_NET_108, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22024(__A22_1__DKCTR1_n, __A22_1__DKCTR2_n, __A22_1__DKCTR1, __A22_1__DKCTR2, __A22_1__DKCTR3_n, __A22_NET_96, GND, __A22_NET_100, __A22_1__DKCTR1_n, __A22_1__DKCTR2, __A22_1__DKCTR3_n, __A22_NET_102, __A22_1__DKCTR3, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22025(__A22_1__DKCTR1, __A22_1__DKCTR2_n, __A22_1__DKCTR1_n, __A22_1__DKCTR2_n, __A22_1__DKCTR3_n, __A22_NET_108, GND, __A22_NET_86, __A22_1__LOW0_n, __A22_NET_91, __A22_1__HIGH0_n, __A22_NET_107, __A22_1__DKCTR3_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22026(__A22_NET_105, WCH34_n, CHWL14_n, __A22_NET_92, __A22_NET_105, __A22_NET_90, GND, __A22_NET_92, CCH34, __A22_NET_90, __A22_1__DATA_n, __A22_1__WDORDR, __A22_NET_95, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22027(__A22_1__HIGH0_n, __A22_NET_92, __A22_1__WRD1BP, __A22_1__WRD1B1, __A22_1__WRD2B2, __A22_NET_87, GND, __A22_NET_88, __A22_1__WRD2B3, __A22_NET_86, __A22_NET_89, __A22_NET_89, __A22_1__LOW1_n, p4VDC, SIM_RST, SIM_CLK);
    U74LVC07 U22028(__A22_NET_87, __A22_1__DATA_n_U22028_2, __A22_NET_88, __A22_1__DATA_n_U22028_4, __A22_NET_229, __A22_1__DATA_n_U22028_6, GND, __A22_1__DATA_n_U22028_8, __A22_NET_274, __A22_1__DATA_n_U22028_10, __A22_NET_263, __A22_1__DATA_n_U22028_12, __A22_NET_187, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22029(__A22_1__DKDAT_n, __A22_NET_95, __A22_1__ORDRBT, __A22_NET_245, WCH34_n, PC15_n, GND, __A22_NET_245, __A22_NET_243, __A22_NET_244, __A22_NET_244, CCH34, __A22_NET_243, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22130(__A22_1__BSYNC_n, __A22_1__RDOUT_n,  ,  ,  ,  , GND,  ,  ,  ,  , DKDATA, __A22_1__DKDAT_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U22131(DKBSNC, __A22_1__BSYNC_n,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22032(__A22_NET_242, WCH34_n, CHWL01_n, __A22_NET_240, __A22_NET_242, __A22_NET_241, GND, __A22_NET_240, CCH34, __A22_NET_241, WCH34_n, CHWL02_n, __A22_NET_252, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22033(__A22_1__HIGH1_n, __A22_NET_240, __A22_1__HIGH1_n, __A22_NET_253, __A22_1__LOW5_n, __A22_NET_230, GND, __A22_NET_231, __A22_1__HIGH0_n, __A22_NET_247, __A22_1__LOW2_n, __A22_1__WRD1B1, __A22_1__LOW6_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22034(__A22_NET_253, __A22_NET_252, __A22_NET_251, __A22_NET_251, __A22_NET_253, CCH34, GND, WCH34_n, CHWL13_n, __A22_NET_246, __A22_NET_246, __A22_NET_248, __A22_NET_247, p4VDC, SIM_RST, SIM_CLK);
    U74HC4002 U22035(__A22_NET_229, __A22_NET_230, __A22_NET_231, __A22_NET_225, __A22_NET_239,  , GND,  , __A22_NET_275, __A22_NET_235, __A22_NET_270, __A22_NET_273, __A22_NET_274, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22036(__A22_NET_248, __A22_NET_247, CCH34, __A22_NET_227, WCH34_n, CHWL12_n, GND, __A22_NET_227, __A22_NET_228, __A22_NET_226, __A22_NET_226, CCH34, __A22_NET_228, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22037(__A22_1__HIGH0_n, __A22_NET_226, __A22_1__HIGH0_n, __A22_NET_222, __A22_1__LOW4_n, __A22_NET_239, GND, __A22_NET_275, __A22_1__HIGH0_n, __A22_NET_236, __A22_1__LOW5_n, __A22_NET_225, __A22_1__LOW3_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22038(__A22_NET_223, WCH34_n, CHWL11_n, __A22_NET_222, __A22_NET_223, __A22_NET_224, GND, __A22_NET_222, CCH34, __A22_NET_224, WCH34_n, CHWL10_n, __A22_NET_237, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22039(__A22_NET_236, __A22_NET_237, __A22_NET_238, __A22_NET_238, __A22_NET_236, CCH34, GND, WCH34_n, CHWL09_n, __A22_NET_232, __A22_NET_232, __A22_NET_234, __A22_NET_233, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22040(__A22_NET_234, __A22_NET_233, CCH34, __A22_NET_276, WCH34_n, CHWL08_n, GND, __A22_NET_276, __A22_NET_280, __A22_NET_279, __A22_NET_279, CCH34, __A22_NET_280, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22041(__A22_1__HIGH0_n, __A22_NET_233, __A22_1__HIGH0_n, __A22_NET_279, __A22_1__LOW7_n, __A22_NET_270, GND, __A22_NET_273, __A22_1__HIGH1_n, __A22_NET_284, __A22_1__LOW0_n, __A22_NET_235, __A22_1__LOW6_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22042(__A22_NET_271, WCH34_n, CHWL07_n, __A22_NET_284, __A22_NET_271, __A22_NET_272, GND, __A22_NET_284, CCH34, __A22_NET_272, WCH34_n, CHWL06_n, __A22_NET_287, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22043(__A22_NET_285, __A22_NET_287, __A22_NET_286, __A22_NET_286, __A22_NET_285, CCH34, GND, WCH34_n, CHWL05_n, __A22_NET_281, __A22_NET_281, __A22_NET_282, __A22_NET_283, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22044(__A22_1__HIGH1_n, __A22_NET_285, __A22_1__HIGH1_n, __A22_NET_283, __A22_1__LOW2_n, __A22_NET_265, GND, __A22_NET_259, __A22_1__HIGH1_n, __A22_NET_254, __A22_1__LOW3_n, __A22_NET_262, __A22_1__LOW1_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22045(__A22_NET_282, __A22_NET_283, CCH34, __A22_NET_266, WCH34_n, CHWL04_n, GND, __A22_NET_266, __A22_NET_255, __A22_NET_254, __A22_NET_254, CCH34, __A22_NET_255, p4VDC, SIM_RST, SIM_CLK);
    U74HC4002 U22046(__A22_NET_263, __A22_NET_262, __A22_NET_265, __A22_NET_259, __A22_NET_261,  , GND,  , __A22_NET_177, __A22_NET_183, __A22_NET_160, __A22_NET_156, __A22_NET_187, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22047(__A22_NET_256, WCH34_n, CHWL03_n, __A22_NET_257, __A22_NET_256, __A22_NET_258, GND, __A22_NET_257, CCH34, __A22_NET_258, WCH35_n, CHWL16_n, __A22_NET_267, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22048(__A22_1__HIGH1_n, __A22_NET_257, __A22_1__HIGH2_n, __A22_NET_269, __A22_1__LOW0_n, __A22_NET_177, GND, __A22_NET_183, __A22_1__HIGH2_n, __A22_NET_180, __A22_1__LOW1_n, __A22_NET_261, __A22_1__LOW4_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22049(__A22_NET_269, __A22_NET_267, __A22_NET_268, __A22_NET_268, __A22_NET_269, CCH35, GND, WCH35_n, CHWL14_n, __A22_NET_182, __A22_NET_182, __A22_NET_181, __A22_NET_180, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22050(__A22_NET_181, __A22_NET_180, CCH35, __A22_NET_176, WCH35_n, CHWL13_n, GND, __A22_NET_176, __A22_NET_175, __A22_NET_174, __A22_NET_174, CCH35, __A22_NET_175, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22051(__A22_1__HIGH2_n, __A22_NET_174, __A22_1__HIGH2_n, __A22_NET_190, __A22_1__LOW3_n, __A22_NET_156, GND, __A22_NET_164, __A22_1__HIGH2_n, __A22_NET_184, __A22_1__LOW4_n, __A22_NET_160, __A22_1__LOW2_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22052(__A22_NET_188, WCH35_n, CHWL12_n, __A22_NET_190, __A22_NET_188, __A22_NET_189, GND, __A22_NET_190, CCH35, __A22_NET_189, WCH35_n, CHWL11_n, __A22_NET_185, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22053(__A22_NET_184, __A22_NET_185, __A22_NET_186, __A22_NET_186, __A22_NET_184, CCH35, GND, WCH35_n, CHWL10_n, __A22_NET_157, __A22_NET_157, __A22_NET_159, __A22_NET_158, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22054(__A22_NET_159, __A22_NET_158, CCH35, __A22_NET_154, WCH35_n, CHWL09_n, GND, __A22_NET_154, __A22_NET_155, __A22_NET_153, __A22_NET_153, CCH35, __A22_NET_155, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22055(__A22_1__HIGH2_n, __A22_NET_158, __A22_1__HIGH2_n, __A22_NET_153, __A22_1__LOW6_n, __A22_NET_168, GND, __A22_NET_167, __A22_1__HIGH2_n, __A22_NET_173, __A22_1__LOW7_n, __A22_NET_161, __A22_1__LOW5_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC4002 U22056(__A22_NET_163, __A22_NET_164, __A22_NET_161, __A22_NET_168, __A22_NET_167,  , GND,  , __A22_NET_215, __A22_NET_214, __A22_NET_195, __A22_NET_194, __A22_NET_213, p4VDC, SIM_RST, SIM_CLK);
    U74LVC07 U22057(__A22_NET_163, __A22_1__DATA_n_U22057_2, __A22_NET_213, __A22_1__DATA_n_U22057_4, __A22_NET_202, __A22_1__DATA_n_U22057_6, GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22058(__A22_NET_172, WCH35_n, CHWL08_n, __A22_NET_173, __A22_NET_172, __A22_NET_171, GND, __A22_NET_173, CCH35, __A22_NET_171, WCH35_n, CHWL07_n, __A22_NET_162, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22059(__A22_NET_170, __A22_NET_162, __A22_NET_169, __A22_NET_169, __A22_NET_170, CCH35, GND, WCH35_n, CHWL06_n, __A22_NET_209, __A22_NET_209, __A22_NET_210, __A22_NET_211, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22060(__A22_1__HIGH3_n, __A22_NET_170, __A22_1__HIGH3_n, __A22_NET_211, __A22_1__LOW1_n, __A22_NET_214, GND, __A22_NET_195, __A22_1__HIGH3_n, __A22_NET_208, __A22_1__LOW2_n, __A22_NET_215, __A22_1__LOW0_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22061(__A22_NET_210, __A22_NET_211, CCH35, __A22_NET_207, WCH35_n, CHWL05_n, GND, __A22_NET_207, __A22_NET_206, __A22_NET_208, __A22_NET_208, CCH35, __A22_NET_206, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22062(__A22_NET_219, WCH35_n, CHWL04_n, __A22_NET_221, __A22_NET_219, __A22_NET_220, GND, __A22_NET_221, CCH35, __A22_NET_220, WCH35_n, CHWL03_n, __A22_NET_217, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22063(__A22_1__HIGH3_n, __A22_NET_221, __A22_1__HIGH3_n, __A22_NET_196, __A22_1__LOW4_n, __A22_1__WRD2B3, GND, __A22_1__WRD2B2, __A22_1__HIGH3_n, __A22_NET_191, __A22_1__LOW5_n, __A22_NET_194, __A22_1__LOW3_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U22064(__A22_NET_196, __A22_NET_217, __A22_NET_218, __A22_NET_218, __A22_NET_196, CCH35, GND, WCH35_n, CHWL02_n, __A22_NET_198, __A22_NET_198, __A22_NET_197, __A22_NET_191, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U22065(__A22_NET_197, __A22_NET_191, CCH35, __A22_NET_192, WCH35_n, CHWL01_n, GND, __A22_NET_192, __A22_NET_204, __A22_NET_203, __A22_NET_203, CCH35, __A22_NET_204, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22066(__A22_1__HIGH3_n, __A22_NET_203, __A22_1__HIGH3_n, __A22_NET_199, __A22_1__LOW7_n, __A22_NET_201, GND,  ,  ,  ,  , __A22_NET_193, __A22_1__LOW6_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U22067(__A22_NET_205, WCH35_n, PC15_n, __A22_NET_199, __A22_NET_205, __A22_NET_200, GND, __A22_NET_199, CCH35, __A22_NET_200, __A22_NET_193, __A22_NET_201, __A22_NET_202, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U22068(__A22_1__BSYNC_n, __A22_1__RDOUT_n, __A22_1__HIGH1_n, __A22_NET_244, __A22_1__LOW7_n, __A22_1__WRD1BP, GND,  ,  ,  ,  , __A22_1__DKDATB, __A22_1__DKDAT_n, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b1, 1'b1) U23001(__A23_1__NOXP, __A23_1__NOXM, __A23_1__NOYM, __A23_1__NOZP, __A23_1__NOZM, __A23_NET_178, GND, __A23_NET_184, __A23_1__MISSX, __A23_1__MISSY, __A23_1__MISSZ, __A23_NET_179, __A23_1__NOYP, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U23002(__A23_NET_179, __A23_NET_185_U23002_2, __A23_NET_178, __A23_NET_185_U23002_4, __A23_NET_175, __A23_NET_174_U23002_6, GND, __A23_NET_174_U23002_8, __A23_NET_173,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1) U23003(F18B, __A23_1__F18B_n, __A23_1__PIPGXp, __A23_NET_208, __A23_1__PIPGXm, __A23_NET_171, GND, __A23_NET_160, F5ASB2, __A23_NET_127, __A23_1__PIPGYp, __A23_NET_126, __A23_1__PIPGYm, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23004(__A23_NET_182, __A23_1__F18B_n, __A23_NET_185, __A23_NET_176, F5ASB0_n, __A23_NET_184, GND, __A23_NET_174, CCH33, PIPAFL, __A23_NET_172, __A23_NET_161, __A23_NET_159, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b1, 1'b0) U23005(__A23_1__BOTHX, __A23_1__BOTHY, __A23_NET_182, __A23_NET_176, PIPAFL, __A23_NET_173, GND, __A23_NET_162, __A23_NET_209, __A23_NET_170, __A23_NET_208, __A23_NET_175, __A23_1__BOTHZ, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23006(__A23_NET_171, __A23_NET_170, PIPPLS_n, SB2_n, __A23_1__P04A, __A23_1__PIPSAM, GND,  ,  ,  ,  , __A23_NET_172, __A23_NET_163, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23007(__A23_NET_161, __A23_NET_159, __A23_NET_162, __A23_NET_164, __A23_NET_160, __A23_NET_159, GND, __A23_NET_161, __A23_NET_160, __A23_NET_165, __A23_NET_164, __A23_NET_163, __A23_NET_209, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23008(__A23_NET_163, __A23_NET_209, __A23_NET_165, __A23_NET_154, __A23_NET_160, __A23_NET_155, GND, __A23_NET_156, __A23_NET_160, __A23_NET_157, __A23_NET_154, __A23_NET_170, __A23_NET_158, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23009(__A23_NET_163, __A23_NET_170, __A23_NET_209, __A23_NET_170, __A23_NET_171, __A23_NET_169, GND, __A23_NET_166, __A23_NET_163, __A23_NET_158, __A23_NET_171, __A23_NET_168, __A23_NET_208, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U23010(__A23_NET_209, __A23_NET_158, __A23_NET_168, __A23_NET_169, __A23_NET_156, __A23_NET_155, GND, __A23_NET_156, __A23_NET_155, __A23_NET_166, __A23_NET_167, __A23_NET_167, __A23_NET_208, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U23011(__A23_NET_170, __A23_NET_158, __A23_NET_157, __A23_1__BOTHX, __A23_NET_171, __A23_NET_208, GND, __A23_1__PIPGXm, __A23_NET_206, __A23_1__NOXM, __A23_1__NOXM, __A23_1__F18AX, __A23_NET_206, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23012(__A23_1__NOXP, __A23_1__PIPGXp, __A23_NET_205, __A23_NET_205, __A23_1__NOXP, __A23_1__F18AX, GND, __A23_1__MISSX, F5ASB2, __A23_NET_211, __A23_NET_126, __A23_NET_127, __A23_1__BOTHY, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b1, 1'b0, 1'b0) U23013(__A23_1__PIPGXp, __A23_1__PIPGXm, __A23_NET_163, __A23_NET_158, __A23_NET_208, PIPXP, GND, PIPXM, __A23_NET_209, __A23_NET_158, __A23_NET_171, __A23_1__MISSX, __A23_NET_211, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23014(__A23_NET_126, __A23_NET_194, __A23_NET_188, __A23_NET_194, __A23_NET_127, __A23_NET_196, GND, __A23_NET_199, __A23_NET_190, __A23_NET_194, __A23_NET_127, __A23_NET_192, __A23_NET_190, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23015(__A23_NET_188, __A23_NET_194, __A23_NET_190, __A23_NET_204, __A23_NET_126, __A23_NET_201, GND, __A23_NET_200, __A23_NET_188, __A23_NET_204, __A23_NET_127, __A23_NET_198, __A23_NET_126, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23016(__A23_NET_193, __A23_NET_192, __A23_NET_195, __A23_NET_195, __A23_NET_193, __A23_NET_196, GND, __A23_NET_189, __A23_NET_193, __A23_NET_109, __A23_NET_195, __A23_NET_189, __A23_NET_187, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b1) U23017(__A23_NET_199, __A23_NET_198, __A23_NET_202, __A23_NET_201, __A23_NET_200, __A23_NET_197, GND, __A23_1__MISSY, __A23_1__PIPGYp, __A23_1__PIPGYm, __A23_NET_129, __A23_NET_202, __A23_NET_197, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0) U23018(F5ASB2, __A23_NET_189, __A23_1__PIPGZp, __A23_NET_143, __A23_1__PIPGZm, __A23_NET_101, GND, __A23_NET_116, F5ASB2, __A23_1__F18A_n, F18A, __A23_1__F18AX, __A23_1__F18A_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U23019(__A23_NET_191, __A23_NET_189, __A23_NET_202, __A23_NET_203, __A23_NET_197, __A23_NET_189, GND, __A23_NET_109, __A23_NET_190, __A23_NET_188, __A23_NET_188, __A23_NET_187, __A23_NET_190, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U23020(__A23_NET_204, __A23_NET_191, __A23_NET_194, __A23_NET_194, __A23_NET_204, __A23_NET_203, GND, __A23_1__PIPGYm, __A23_NET_120, __A23_1__NOYM, __A23_1__NOYM, __A23_1__F18AX, __A23_NET_120, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23021(__A23_1__NOYP, __A23_1__PIPGYp, __A23_NET_123, __A23_NET_123, __A23_1__NOYP, __A23_1__F18AX, GND, __A23_1__MISSY, F5ASB2, __A23_NET_129, __A23_NET_101, __A23_NET_143, __A23_1__BOTHZ, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23022(__A23_NET_190, __A23_NET_204, __A23_NET_188, __A23_NET_204, __A23_NET_126, PIPYM, GND, __A23_NET_105, __A23_NET_101, __A23_NET_148, __A23_NET_107, PIPYP, __A23_NET_127, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23023(__A23_NET_108, __A23_NET_148, __A23_NET_107, __A23_NET_148, __A23_NET_143, __A23_NET_119, GND, __A23_NET_118, __A23_NET_108, __A23_NET_148, __A23_NET_101, __A23_NET_104, __A23_NET_143, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b0, 1'b1) U23024(__A23_NET_107, __A23_NET_111, __A23_NET_108, __A23_NET_111, __A23_NET_143, __A23_NET_147, GND, __A23_1__MISSZ, __A23_1__PIPGZp, __A23_1__PIPGZm, __A23_NET_149, __A23_NET_115, __A23_NET_101, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U23025(__A23_NET_102, __A23_NET_105, __A23_NET_103, __A23_NET_103, __A23_NET_102, __A23_NET_104, GND, __A23_1__PIPGZm, __A23_NET_144, __A23_1__NOZM, __A23_1__NOZM, __A23_1__F18AX, __A23_NET_144, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 #(1'b0, 1'b1, 1'b0) U23026(__A23_NET_119, __A23_NET_118, __A23_NET_112, __A23_NET_115, __A23_NET_147, __A23_NET_117, GND, PIPZP, __A23_NET_107, __A23_NET_111, __A23_NET_143, __A23_NET_112, __A23_NET_117, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23027(__A23_1__NOZP, __A23_1__PIPGZp, __A23_NET_153, __A23_NET_153, __A23_1__NOZP, __A23_1__F18AX, GND, __A23_1__MISSZ, F5ASB2, __A23_NET_149, __A23_NET_116, __A23_NET_102, __A23_NET_110, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23028(__A23_NET_106, __A23_NET_103, __A23_NET_116, __A23_NET_113, __A23_NET_116, __A23_NET_112, GND, __A23_NET_117, __A23_NET_116, __A23_NET_114, __A23_NET_110, __A23_NET_107, __A23_NET_108, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U23029(__A23_NET_107, __A23_NET_108, __A23_NET_106, __A23_NET_111, __A23_NET_113, __A23_NET_148, GND, __A23_NET_111, __A23_NET_114, __A23_NET_148, CHWL16_n, WCH14_n, __A23_NET_252, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23030(__A23_NET_108, __A23_NET_111, __A23_NET_250, CCH14, __A23_NET_257, __A23_NET_253, GND, __A23_NET_255, __A23_NET_245, CCH14, __A23_NET_244, PIPZM, __A23_NET_101, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23031(__A23_NET_250, __A23_NET_252, __A23_NET_253, CH1416, RCH14_n, __A23_NET_250, GND, __A23_NET_250, F5ASB2_n, CDUXD, XB0_n, __A23_NET_268, __A23_NET_251, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0) U23032(__A23_NET_251, __A23_NET_256, OCTAD5, __A23_NET_268, __A23_NET_246, __A23_NET_243, GND, __A23_NET_267, __A23_NET_266, __A23_NET_270, __A23_NET_269, __A23_NET_264, __A23_NET_263, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23033(CDUXDP, POUT_n, __A23_NET_256, CDUXDM, MOUT_n, __A23_NET_256, GND, ZOUT_n, __A23_NET_256, __A23_NET_257, CHWL14_n, WCH14_n, __A23_NET_254, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23034(__A23_NET_245, __A23_NET_254, __A23_NET_255, CH1414, RCH14_n, __A23_NET_245, GND, __A23_NET_245, F5ASB2_n, CDUYD, XB1_n, __A23_NET_268, __A23_NET_246, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23035(CDUYDP, POUT_n, __A23_NET_243, CDUYDM, MOUT_n, __A23_NET_243, GND, ZOUT_n, __A23_NET_243, __A23_NET_244, CHWL13_n, WCH14_n, __A23_NET_249, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23036(__A23_NET_248, __A23_NET_249, __A23_NET_247, CH1413, RCH14_n, __A23_NET_248, GND, __A23_NET_248, F5ASB2_n, CDUZD, XB2_n, __A23_NET_268, __A23_NET_266, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23037(__A23_NET_248, CCH14, __A23_NET_273, CCH14, __A23_NET_260, __A23_NET_272, GND, __A23_NET_259, __A23_NET_261, CCH14, __A23_NET_262, __A23_NET_247, __A23_NET_265, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23038(CDUZDP, POUT_n, __A23_NET_267, CDUZDM, MOUT_n, __A23_NET_267, GND, ZOUT_n, __A23_NET_267, __A23_NET_265, CHWL12_n, WCH14_n, __A23_NET_271, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23039(__A23_NET_273, __A23_NET_271, __A23_NET_272, CH1412, RCH14_n, __A23_NET_273, GND, __A23_NET_273, F5ASB2_n, TRUND, XB3_n, __A23_NET_268, __A23_NET_269, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23040(TRNDP, POUT_n, __A23_NET_270, TRNDM, MOUT_n, __A23_NET_270, GND, ZOUT_n, __A23_NET_270, __A23_NET_260, CHWL11_n, WCH14_n, __A23_NET_258, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23041(__A23_NET_261, __A23_NET_258, __A23_NET_259, CH1411, RCH14_n, __A23_NET_261, GND, __A23_NET_261, F5ASB2_n, SHAFTD, XB4_n, __A23_NET_268, __A23_NET_263, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23042(SHFTDP, POUT_n, __A23_NET_264, SHFTDM, MOUT_n, __A23_NET_264, GND, ZOUT_n, __A23_NET_264, __A23_NET_262, CHWL05_n, __A23_2__WCH07_n, __A23_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23043(__A23_NET_219, __A23_NET_222, E5, E5, __A23_NET_219, __A23_2__CCH07, GND, __A23_2__RCH07_n, __A23_NET_219, CH0705, CHWL06_n, __A23_2__WCH07_n, __A23_NET_220, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23044(__A23_NET_223, __A23_NET_220, E6, E6, __A23_NET_223, __A23_2__CCH07, GND, __A23_2__RCH07_n, __A23_NET_223, CH0706, CHWL07_n, __A23_2__WCH07_n, __A23_NET_227, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23045(E7_n, __A23_NET_227, __A23_NET_225, __A23_NET_225, E7_n, __A23_2__CCH07, GND, __A23_2__RCH07_n, E7_n, CH0707, XB7_n, XT0_n, __A23_NET_212, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U23046(WCHG_n, XT0_n, CCHG_n, XB7_n, XT0_n, __A23_2__CCH07, GND, __A23_NET_229, T6ON_n, T6RPT, CCH13, __A23_NET_214, XB7_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U23047(__A23_NET_214, __A23_2__WCH07_n, __A23_NET_212, __A23_2__RCH07_n, __A23_NET_218, __A23_2__OT1108, GND, __A23_2__OT1113, __A23_NET_238, __A23_2__OT1114, __A23_NET_237, __A23_2__OT1116, __A23_NET_242, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23048(__A23_NET_213, CHWL08_n, WCH11_n, __A23_NET_218, __A23_NET_213, __A23_NET_217, GND, __A23_NET_218, CCH11, __A23_NET_217, RCH11_n, __A23_NET_218, CH1108, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23049(__A23_NET_216, CHWL13_n, WCH11_n, __A23_NET_238, __A23_NET_216, __A23_NET_215, GND, __A23_NET_238, CCH11, __A23_NET_215, RCH11_n, __A23_NET_238, CH1113, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23050(__A23_NET_236, CHWL14_n, WCH11_n, __A23_NET_237, __A23_NET_236, __A23_NET_235, GND, __A23_NET_237, CCH11, __A23_NET_235, RCH11_n, __A23_NET_237, CH1114, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23051(__A23_NET_241, CHWL16_n, WCH11_n, __A23_NET_242, __A23_NET_241, __A23_NET_240, GND, __A23_NET_242, CCH11, __A23_NET_240, RCH11_n, __A23_NET_242, CH1116, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23052(__A23_NET_231, CHWL16_n, WCH12_n, __A23_NET_230, __A23_NET_231, __A23_NET_239, GND, __A23_NET_230, CCH12, __A23_NET_239, RCH12_n, __A23_NET_230, CH1216, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0) U23053(__A23_NET_230, __A23_2__ISSTDC,  ,  , __A23_NET_232, ALTEST, GND, __A23_1__P04A, P04_n, __A23_1__PIPSAM_n, __A23_1__PIPSAM, __A23_1__PIPAXp_n, PIPAXp, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U23054(__A23_NET_228, CHWL16_n, WCH13_n, T6ON_n, __A23_NET_228, __A23_NET_229, GND, RCH13_n, T6ON_n, CH1316, CHWL10_n, WCH13_n, __A23_NET_234, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b0) U23055(__A23_NET_232, __A23_NET_234, __A23_NET_233, __A23_NET_233, __A23_NET_232, CCH13, GND, RCH13_n, __A23_NET_232, CH1310, __A23_1__PIPSAM_n, __A23_1__PIPAXp_n, __A23_1__PIPGXp, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U23056(PIPAXm, __A23_1__PIPAXm_n, PIPAYp, __A23_1__PIPAYp_n, PIPAYm, __A23_1__PIPAYm_n, GND, __A23_1__PIPAZp_n, PIPAZp, __A23_1__PIPAZm_n, PIPAZm,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23057(__A23_1__PIPGXm, __A23_1__PIPSAM_n, __A23_1__PIPAXm_n, __A23_1__PIPGYp, __A23_1__PIPSAM_n, __A23_1__PIPAYp_n, GND, __A23_1__PIPSAM_n, __A23_1__PIPAYm_n, __A23_1__PIPGYm, __A23_1__PIPSAM_n, __A23_1__PIPAZp_n, __A23_1__PIPGZp, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U23058(__A23_1__PIPGZm, __A23_1__PIPSAM_n, __A23_1__PIPAZm_n,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U24001(WL01, CHWL01_n, WL02, CHWL02_n, WL03, CHWL03_n, GND, CHWL04_n, WL04, CHWL05_n, WL05, CHWL06_n, WL06, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U24002(WL07, CHWL07_n, WL08, CHWL08_n, WL09, CHWL09_n, GND, CHWL10_n, WL10, CHWL11_n, WL11, CHWL12_n, WL12, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U24003(WL13, CHWL13_n, WL14, CHWL14_n, WL16, CHWL16_n, GND, RCHAT_n, __A24_NET_212, RCHBT_n, __A24_NET_213,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U24104(PIPASW, PIPPLS_n, SB1_n, PIPDAT, PIPPLS_n, SB2_n, GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U24105(FS04, __A24_NET_217, F03B, __A24_1__F03B_n, __A24_NET_220, PIPPLS_n, GND,  ,  ,  ,  ,  ,  , p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U24106(__A24_1__F03B_n, __A24_NET_217, FS05, SB0_n, __A24_NET_216, __A24_1__3200C, GND, __A24_1__3200D, __A24_NET_216, SB0_n, FS05_n, __A24_NET_220, FS05, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U24107(__A24_1__PIPINT, PIPPLS_n, __A24_NET_215, __A24_1__800SET, __A24_1__F07A_n, SB1_n, GND, F07B_n, SB1_n, __A24_1__800RST, F05A_n, SB0_n, __A24_1__3200A, p4VDC, SIM_RST, SIM_CLK);
    U74HC04 U24108(SB4, __A24_NET_215, F07A, __A24_1__F07A_n, F04B, __A24_NET_216, GND, __A24_NET_202, F02B, __A24_NET_201, F01B, __A24_NET_203, F01A, p4VDC, SIM_RST, SIM_CLK);
    U74HC02 U24109(__A24_1__3200B, F05B_n, SB0_n, __A24_1__CDUCLK, __A24_NET_203, SB0_n, GND, F05B_n, SB1_n, __A24_1__RRRST, F05B_n, SB1_n, __A24_1__LRRST, p4VDC, SIM_RST, SIM_CLK);
    U74HC27 U24110(FS03, __A24_NET_202, SB0_n, FS02, __A24_NET_201, __A24_1__25KPPS, GND,  ,  ,  ,  , __A24_1__12KPPS, SB0_n, p4VDC, SIM_RST, SIM_CLK);
    U74LVC07 U24011(__A24_NET_247, CHOR01_n_U24011_2, __A24_NET_246, CHOR02_n_U24011_4, __A24_NET_248, CHOR03_n_U24011_6, GND, CHOR04_n_U24011_8, __A24_NET_241, CHOR05_n_U24011_10, __A24_NET_245, CHOR06_n_U24011_12, __A24_NET_244, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U24012(CH01, CHOR01_n, RCHG_n, CH02, CHOR02_n, RCHG_n, GND, CHOR03_n, RCHG_n, CH03, CHOR04_n, RCHG_n, CH04, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U24013(CHAT02, CHBT02, CHAT03, CHBT03, CH1603, __A24_NET_248, GND, __A24_NET_241, CHAT04, CHBT04, CH1604, __A24_NET_246, CH1602, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U24014(CH05, CHOR05_n, RCHG_n, CH06, CHOR06_n, RCHG_n, GND, CHOR07_n, RCHG_n, CH07, CHOR08_n, RCHG_n, CH08, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U24015(__A24_NET_245, CHAT05, CHBT05, CH1605, CH1505,  , GND,  , CHAT08, CHBT08, CH1108, CH1208, __A24_NET_256, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U24016(CHAT06, CHBT06, CHAT07, CHBT07, CH1607, __A24_NET_253, GND, __A24_NET_250, CH1109, CH1209, CH3209, __A24_NET_244, CH1606, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U24017(__A24_NET_253, CHOR07_n_U24017_2, __A24_NET_256, CHOR08_n_U24017_4, __A24_NET_249, CHOR09_n_U24017_6, GND, CHOR09_n_U24017_8, __A24_NET_250, CHOR10_n_U24017_10, __A24_NET_251, CHOR10_n_U24017_12, __A24_NET_252, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U24018(CH09, CHOR09_n, RCHG_n, __A24_NET_249, CHAT09, CHBT09, GND, CHOR10_n, RCHG_n, CH10, CHAT10, CHBT10, __A24_NET_251, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U24019(CH1110, CH1210, CH1111, CH1211, CH3311, __A24_NET_229, GND, __A24_NET_226, CH1116, CH1216, CH3316, __A24_NET_252, CH3210, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U24020(CH11, CHOR11_n, RCHG_n, __A24_NET_228, CHAT11, CHBT11, GND, CHOR12_n, RCHG_n, CH12, CHOR13_n, RCHG_n, CH13, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U24021(__A24_NET_228, CHOR11_n_U24021_2, __A24_NET_229, CHOR11_n_U24021_4, __A24_NET_230, CHOR12_n_U24021_6, GND, CHOR13_n_U24021_8, __A24_NET_222, CHOR14_n_U24021_10, __A24_NET_223, CHOR16_n_U24021_12, __A24_NET_226, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U24022(__A24_NET_230, CHAT12, CHBT12, CH1112, CH1212,  , GND,  , CHAT13, CHBT13, CH1113, CH3313, __A24_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b0, 1'b1) U24023(CH14, CHOR14_n, RCHG_n, CH16, CHOR16_n, RCHG_n, GND, T08, CDUSTB_n, __A24_NET_238, __A24_NET_238, T06, CDUSTB_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U24024(__A24_NET_223, CHAT14, CHBT14, CH1114, CH3314,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U24025(FLASH, FS17, FS16, __A24_NET_234, FS08, FS09, GND, __A24_NET_195, GOJAM, __A24_NET_196, __A24_NET_200, GOJAM, __A24_NET_199, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U24026(FLASH, FLASH_n, __A24_NET_239, __A24_NET_240, GTSET, GTSET_n, GND, GTRST_n, __A24_NET_235, __A24_2__FS06_n, FS06, __A24_2__FS08_n, FS08, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U24027(FS07_n, __A24_2__FS08_n, __A24_2__FS06_n, F05B_n, __A24_NET_240, GTSET, GND, __A24_NET_235, __A24_NET_240, F05B_n, FS06, __A24_NET_239, FS09_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U24028(FS06, F05B_n, CCHG_n, XT1_n, XB3_n, __A24_NET_195, GND, __A24_NET_205, WCHG_n, XT1_n, XB3_n, __A24_NET_233, FS07A, p4VSW, SIM_RST, SIM_CLK);
    U74LVC07 U24029(__A24_NET_233, GTONE_U24029_2, __A24_NET_234, GTONE_U24029_4,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U24030(__A24_NET_196, CCH13, __A24_NET_199, CCH14, __A24_NET_197, CCH34, GND, CCH35, __A24_NET_208, RCH13_n, __A24_NET_211, RCH14_n, __A24_NET_210, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U24031(CCHG_n, XT1_n, CCHG_n, XT3_n, XB4_n, __A24_NET_198, GND, __A24_NET_209, CCHG_n, XT3_n, XB5_n, __A24_NET_200, XB4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U24032(__A24_NET_197, __A24_NET_198, GOJAM, __A24_NET_208, __A24_NET_209, GOJAM, GND, XT1_n, XB3_n, __A24_NET_211, XT1_n, XB4_n, __A24_NET_210, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0) U24033(__A24_NET_205, WCH13_n, __A24_NET_204, WCH14_n, __A24_NET_207, WCH34_n, GND, WCH35_n, __A24_NET_206,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U24034(WCHG_n, XT1_n, WCHG_n, XT3_n, XB4_n, __A24_NET_207, GND, __A24_NET_206, WCHG_n, XT3_n, XB5_n, __A24_NET_204, XB4_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U24035(__A24_NET_212, XB4_n, XT0_n, __A24_NET_213, XT0_n, XB3_n, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U24036(FS07A, __A24_NET_219, __A24_NET_219, ELSNCN, __A24_NET_219, ELSNCM, GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U24037(CHAT01, CHBT01,  ,  ,  ,  , GND,  ,  ,  ,  , __A24_NET_247, CH1601, p4VSW, SIM_RST, SIM_CLK);
    U74LVC06 U24038(FS07A, MON800_U24038_2,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    SST39VF200A U31001(__B01_1__FADDR16, __B01_1__FADDR15, __B01_1__FADDR14, __B01_1__FADDR13, __B01_1__FADDR12, __B01_1__FADDR11, __B01_1__FADDR10, __B01_1__FADDR9,  ,  , p4VSW,  ,  ,  ,  ,  ,  , __B01_1__FADDR8, __B01_1__FADDR7, __B01_1__FADDR6, __B01_1__FADDR5, __B01_1__FADDR4, __B01_1__FADDR3, __B01_1__FADDR2, __B01_1__FADDR1, __B01_NET_166, GND, __B01_NET_118, SA01_U31001_29, SA09_U31001_30, SA02_U31001_31, SA10_U31001_32, SA03_U31001_33, SA11_U31001_34, SA04_U31001_35, SA12_U31001_36, p4VSW, SA05_U31001_38, SA13_U31001_39, SA06_U31001_40, SA14_U31001_41, SA07_U31001_42, SAP_U31001_43, SA08_U31001_44, SA16_U31001_45, GND,  , GND, SIM_RST, SIM_CLK);
    U74HC04 U31002(ROPER, __B01_NET_180, ROPES, __B01_NET_159, ROPET, __B01_NET_152, GND, __B01_NET_186, STR14, __B01_NET_187, STR58, __B01_NET_179, STR912, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U31003(__B01_NET_152, LOMOD, ROPER, __B01_NET_149, __B01_NET_150, __B01_1__FADDR15, GND, __B01_NET_149, ROPES, LOMOD, STR14, __B01_1__FADDR16, STR14, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U31004(ROPET, HIMOD, ROPER, LOMOD, STR14, __B01_NET_155, GND, __B01_NET_156, ROPET, LOMOD, __B01_NET_186, __B01_NET_150, STR912, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U31005(__B01_NET_158, __B01_NET_159, __B01_NET_179, __B01_NET_157, __B01_NET_180, HIMOD, GND, HIMOD, STR58, __B01_NET_188, LOMOD, __B01_NET_187, __B01_NET_189, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U31006(__B01_1__FADDR14, __B01_NET_158, __B01_NET_155, __B01_NET_156, __B01_NET_157,  , GND,  , __B01_NET_184, __B01_NET_162, __B01_NET_154, __B01_NET_181, __B01_1__FADDR13, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U31007(ROPES, HIMOD, ROPES, LOMOD, STR14, __B01_NET_162, GND, __B01_NET_154, __B01_NET_159, HIMOD, __B01_NET_179, __B01_NET_184, STR912, p4VSW, SIM_RST, SIM_CLK);
    U74HC27 U31008(__B01_NET_159, LOMOD, RSTKX_n, RSTKY_n, ZID, __B01_2__RESETK, GND, __B01_1__NOROPE, ROPER, ROPES, ROPET, __B01_NET_181, __B01_NET_186, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U31009(__B01_1__FADDR12, __B01_NET_188, __B01_NET_189, __B01_1__FADDR11, STR210, STR19, GND, STR19, STR311, __B01_1__FADDR10, __B01_1__QUARTERB, __B01_1__QUARTERA, __B01_1__FADDR9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31010(__B01_1__FADDR8, __B01_1__QUARTERA, __B01_1__QUARTERC, __B01_NET_101, __B01_NET_95, __B01_1__QUARTERA, GND, __B01_NET_101, __B01_1__CQA, __B01_1__QUARTERA, __B01_NET_96, __B01_NET_98, __B01_NET_95, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 U31011(IL07, __B01_1__FADDR7, IL06, __B01_1__FADDR6, IL05, __B01_1__FADDR5, GND, __B01_1__FADDR4, IL04, __B01_1__FADDR3, IL03, __B01_1__FADDR2, IL02, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1) U31012(IL01, __B01_1__FADDR1, __B01_NET_133, __B01_NET_118, SETAB, __B01_NET_96, GND, __B01_NET_98, RESETB, __B01_NET_212, __B01_NET_211, __B01_NET_112, __B01_NET_111, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 #(1'b1, 1'b0) U31013(__B01_NET_166, STR19, STR210, STR311, STR412,  , GND,  , XB1E, XB3E, XB5E, XB7E, __B01_2__ES01_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31014(__B01_NET_109, RESETA, __B01_NET_108, __B01_NET_110, __B01_NET_109, __B01_NET_111, GND, __B01_NET_110, RESETA, __B01_NET_111, __B01_NET_96, __B01_NET_144, __B01_NET_143, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1) U31015(__B01_NET_112, __B01_NET_113, __B01_NET_113, __B01_NET_107, __B01_NET_147, __B01_NET_104, GND, __B01_NET_103, __B01_NET_104, __B01_NET_106, __B01_NET_103, __B01_NET_105, __B01_NET_106, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1) U31016(__B01_NET_107, __B01_NET_108, RESETA, __B01_NET_144, SETCD, __B01_NET_140, GND, __B01_NET_142, RESETD, __B01_1__CQA, __B01_NET_148, __B01_NET_242, ZID, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b1, 1'b0) U31017(__B01_NET_141, __B01_NET_143, __B01_1__QUARTERB, __B01_1__QUARTERB, __B01_NET_141, __B01_1__CQB, GND, __B01_NET_139, __B01_1__QUARTERC, __B01_NET_138, __B01_NET_138, __B01_1__CQC, __B01_1__QUARTERC, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 U31018(__B01_NET_139, __B01_NET_140, __B01_NET_142, __B01_NET_148, CLROPE, __B01_NET_109, GND, YB1E, YB3E, __B01_2__ES07_n, YB2E, YB3E, __B01_2__ES08_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U31019(__B01_2__ES02_n, XB2E, XB3E, XB6E, XB7E,  , GND,  , XB4E, XB5E, XB6E, XB7E, __B01_2__ES03_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U31020(__B01_2__ES04_n, XT1E, XT3E, XT5E, XT7E,  , GND,  , XT2E, XT3E, XT6E, XT7E, __B01_2__ES05_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U31021(__B01_2__ES06_n, XT4E, XT5E, XT6E, XT7E,  , GND,  , YT1E, YT3E, YT5E, YT7E, __B01_2__ES09_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC4002 U31022(__B01_2__ES10_n, YT2E, YT3E, YT6E, YT7E,  , GND,  , YT4E, YT5E, YT6E, YT7E, __B01_2__ES11_n, p4VSW, SIM_RST, SIM_CLK);
    U74HC244 U31023(__B01_NET_242, GEMP, SA07_U31023_3, GEM01, SA06_U31023_5, GEM02, SA05_U31023_7, GEM03, SA04_U31023_9, GND, GEM04, SA03_U31023_12, GEM05, SA02_U31023_14, GEM06, SA01_U31023_16, GEM07, SAP_U31023_18, __B01_NET_242, p4VSW, SIM_RST, SIM_CLK);
    U74HC244 U31024(__B01_NET_242, GEM08, SA16_U31024_3, GEM09, SA14_U31024_5, GEM10, SA13_U31024_7, GEM11, SA12_U31024_9, GND, GEM12, SA11_U31024_12, GEM13, SA10_U31024_14, GEM14, SA09_U31024_16, GEM16, SA08_U31024_18, __B01_NET_242, p4VSW, SIM_RST, SIM_CLK);
    MR0A16A U31025(__B01_2__RADDR1, __B01_2__RADDR2, __B01_2__RADDR3, __B01_2__RADDR4, __B01_2__RADDR5, GND, SA01_U31025_7, SA02_U31025_8, SA03_U31025_9, SA04_U31025_10, p4VSW, GND, SA05_U31025_13, SA06_U31025_14, SA07_U31025_15, SA08_U31025_16, __B01_NET_210, __B01_2__RADDR6, __B01_2__RADDR7, __B01_2__RADDR8, __B01_2__RADDR9, __B01_2__RADDR10, __B01_2__RADDR11, GND, GND, GND, p4VSW,  , SA09_U31025_29, SA10_U31025_30, SA11_U31025_31, SA12_U31025_32, p4VSW, GND, SA13_U31025_35, SA14_U31025_36, SAP_U31025_37, SA16_U31025_38, GND, GND, __B01_NET_204, GND, GND, GND, SIM_RST, SIM_CLK, SA01, SA02, SA03, SA04, SA05, SA06, SA07, SA08, SA09, SA10, SA11, SA12, SA13, SA14, SAP, SA16);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31026(__B01_NET_223, __B01_NET_202, __B01_NET_203, __B01_NET_197, __B01_2__ES01_n, __B01_NET_240, GND, __B01_NET_197, __B01_2__RADDR1, __B01_NET_205, __B01_NET_205, __B01_2__RESETK, __B01_2__RADDR1, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1) U31027(WEX, __B01_NET_202, WEY, __B01_NET_203, __B01_NET_224, __B01_NET_218, GND, __B01_NET_204, SBE, __B01_NET_240, SETEK, __B01_NET_221, __B01_NET_222, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31028(__B01_NET_199, __B01_2__ES02_n, __B01_NET_240, __B01_NET_198, __B01_NET_199, __B01_2__RADDR2, GND, __B01_NET_198, __B01_2__RESETK, __B01_2__RADDR2, __B01_2__ES03_n, __B01_NET_240, __B01_NET_201, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31029(__B01_NET_200, __B01_NET_201, __B01_2__RADDR3, __B01_2__RADDR3, __B01_NET_200, __B01_2__RESETK, GND, __B01_2__ES04_n, __B01_NET_240, __B01_NET_192, __B01_NET_192, __B01_2__RADDR4, __B01_NET_191, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31030(__B01_2__RADDR4, __B01_NET_191, __B01_2__RESETK, __B01_NET_194, __B01_2__ES05_n, __B01_NET_240, GND, __B01_NET_194, __B01_2__RADDR5, __B01_NET_190, __B01_NET_190, __B01_2__RESETK, __B01_2__RADDR5, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31031(__B01_NET_241, __B01_2__ES06_n, __B01_NET_240, __B01_NET_196, __B01_NET_241, __B01_2__RADDR6, GND, __B01_NET_196, __B01_2__RESETK, __B01_2__RADDR6, __B01_2__ES07_n, __B01_NET_240, __B01_NET_236, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31032(__B01_NET_235, __B01_NET_236, __B01_2__RADDR7, __B01_2__RADDR7, __B01_NET_235, __B01_2__RESETK, GND, __B01_2__ES08_n, __B01_NET_240, __B01_NET_239, __B01_NET_239, __B01_2__RADDR8, __B01_NET_238, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31033(__B01_2__RADDR8, __B01_NET_238, __B01_2__RESETK, __B01_NET_226, __B01_2__ES09_n, __B01_NET_240, GND, __B01_NET_226, __B01_2__RADDR9, __B01_NET_225, __B01_NET_225, __B01_2__RESETK, __B01_2__RADDR9, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b0, 1'b0) U31034(__B01_NET_230, __B01_2__ES10_n, __B01_NET_240, __B01_NET_229, __B01_NET_230, __B01_2__RADDR10, GND, __B01_NET_229, __B01_2__RESETK, __B01_2__RADDR10, __B01_2__ES11_n, __B01_NET_240, __B01_NET_233, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b1, 1'b0, 1'b0, 1'b1) U31035(__B01_NET_232, __B01_NET_233, __B01_2__RADDR11, __B01_NET_127, CLROPE, __B01_NET_145, GND, __B01_NET_218, __B01_NET_217, __B01_2__EDESTROY, __B01_2__EDESTROY, __B01_NET_222, __B01_NET_220, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31036(__B01_NET_222, __B01_NET_220, __B01_NET_218, __B01_NET_145, RESETB, __B01_NET_105, GND, __B01_NET_145, __B01_NET_147, __B01_NET_146, __B01_NET_146, RESETB, __B01_NET_147, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1) U31037(__B01_NET_221, __B01_NET_211, __B01_NET_127, __B01_1__CQB, __B01_NET_212, __B01_NET_214, GND, __B01_NET_213, __B01_NET_214, __B01_NET_216, __B01_NET_213, __B01_NET_215, __B01_NET_216, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1) U31038(__B01_NET_215, __B01_NET_217, __B01_NET_136, __B01_1__CQC, __B01_NET_125, __B01_NET_128, GND, __B01_NET_129, __B01_NET_128, __B01_NET_131, __B01_NET_129, __B01_NET_130, __B01_NET_131, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b0, 1'b1, 1'b0) U31039(__B01_NET_136, CLROPE, __B01_NET_124, __B01_NET_124, RESETC, __B01_NET_130, GND, __B01_NET_124, __B01_NET_125, __B01_NET_123, __B01_NET_123, RESETC, __B01_NET_125, p4VSW, SIM_RST, SIM_CLK);
    U74HC02 #(1'b0, 1'b1, 1'b1, 1'b0) U31040(__B01_2__RADDR11, __B01_NET_232, __B01_2__RESETK, __B01_NET_224, REX, REY, GND, __B01_NET_223, __B01_2__EDESTROY, __B01_NET_210, __B01_NET_134, __B01_1__NOROPE, __B01_NET_133, p4VSW, SIM_RST, SIM_CLK);
    U74HC04 #(1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0) U31041(SBF, __B01_NET_134,  ,  ,  ,  , GND,  ,  ,  ,  ,  ,  , p4VSW, SIM_RST, SIM_CLK);
    assign MBR1 = MBR1_U4066_8;
    assign MBR2 = MBR2_U4066_10;
    assign MCTRAL_n = MCTRAL_n_U13051_12;
    assign MGOJAM = MGOJAM_U2148_6;
    assign MIIP = MIIP_U3053_6;
    assign MINHL = MINHL_U3053_4;
    assign MINKL = MINKL_U13053_4;
    assign MNISQ = MNISQ_U5068_2;
    assign MON800 = MON800_U24038_2;
    assign MONWT = MONWT_U2148_2;
    assign MOSCAL_n = MOSCAL_n_U13053_2;
    assign MPAL_n = MPAL_n_U12050_2;
    assign MPIPAL_n = MPIPAL_n_U13052_4;
    assign MRAG = MRAG_U7040_2;
    assign MRCH = MRCH_U6058_2;
    assign MREQIN = MREQIN_U13053_6;
    assign MRGG = MRGG_U7039_12;
    assign MRLG = MRLG_U7040_4;
    assign MRPTAL_n = MRPTAL_n_U13051_8;
    assign MRSC = MRSC_U4067_2;
    assign MRULOG = MRULOG_U7040_6;
    assign MSCAFL_n = MSCAFL_n_U13052_10;
    assign MSCDBL_n = MSCDBL_n_U13052_6;
    assign MSQ10 = MSQ10_U3053_2;
    assign MSQ11 = MSQ11_U3054_12;
    assign MSQ12 = MSQ12_U3054_10;
    assign MSQ13 = MSQ13_U3054_8;
    assign MSQ14 = MSQ14_U3054_6;
    assign MSQ16 = MSQ16_U3054_4;
    assign MSQEXT = MSQEXT_U3054_2;
    assign MST1 = MST1_U4066_2;
    assign MST2 = MST2_U4066_4;
    assign MST3 = MST3_U4066_6;
    assign MSTPIT_n = MSTPIT_n_U2148_8;
    assign MT01 = MT01_U2046_2;
    assign MT02 = MT02_U2046_4;
    assign MT03 = MT03_U2046_6;
    assign MT04 = MT04_U2046_8;
    assign MT05 = MT05_U2046_10;
    assign MT06 = MT06_U2046_12;
    assign MT07 = MT07_U2047_2;
    assign MT08 = MT08_U2047_4;
    assign MT09 = MT09_U2047_6;
    assign MT10 = MT10_U2047_8;
    assign MT11 = MT11_U2047_10;
    assign MT12 = MT12_U2047_12;
    assign MTCAL_n = MTCAL_n_U13051_10;
    assign MTCSA_n = MTCSA_n_U3053_8;
    assign MVFAIL_n = MVFAIL_n_U13052_2;
    assign MWAG = MWAG_U7038_12;
    assign MWARNF_n = MWARNF_n_U13052_12;
    assign MWATCH_n = MWATCH_n_U13052_8;
    assign MWBBEG = MWBBEG_U7039_10;
    assign MWBG = MWBG_U7038_4;
    assign MWCH = MWCH_U4066_12;
    assign MWEBG = MWEBG_U7039_6;
    assign MWFBG = MWFBG_U7039_8;
    assign MWG = MWG_U7038_6;
    assign MWL01 = MWL01_U8068_2;
    assign MWL02 = MWL02_U8068_4;
    assign MWL03 = MWL03_U8068_6;
    assign MWL04 = MWL04_U8068_8;
    assign MWL05 = MWL05_U9068_2;
    assign MWL06 = MWL06_U9068_4;
    assign MWL07 = MWL07_U9068_6;
    assign MWL08 = MWL08_U9068_8;
    assign MWL09 = MWL09_U10068_2;
    assign MWL10 = MWL10_U10068_4;
    assign MWL11 = MWL11_U10068_6;
    assign MWL12 = MWL12_U10068_8;
    assign MWL13 = MWL13_U11068_2;
    assign MWL14 = MWL14_U11068_4;
    assign MWL15 = MWL15_U11068_6;
    assign MWL16 = MWL16_U11068_8;
    assign MWLG = MWLG_U7038_10;
    assign MWQG = MWQG_U7039_4;
    assign MWSG = MWSG_U7039_2;
    assign MWYG = MWYG_U7038_2;
    assign MWZG = MWZG_U7038_8;
    assign A2X_n = A2X_n_U5012_10 & A2X_n_U5044_8 & A2X_n_U6004_6;
    assign CHOR01_n = CHOR01_n_U16004_2 & CHOR01_n_U16021_6 & CHOR01_n_U17003_2 & CHOR01_n_U17027_10 & CHOR01_n_U24011_2;
    assign CHOR02_n = CHOR02_n_U16004_4 & CHOR02_n_U16021_8 & CHOR02_n_U17003_4 & CHOR02_n_U17041_2 & CHOR02_n_U24011_4;
    assign CHOR03_n = CHOR03_n_U16004_6 & CHOR03_n_U16021_10 & CHOR03_n_U17003_6 & CHOR03_n_U17041_4 & CHOR03_n_U24011_6;
    assign CHOR04_n = CHOR04_n_U16004_8 & CHOR04_n_U16021_12 & CHOR04_n_U17003_8 & CHOR04_n_U17041_6 & CHOR04_n_U24011_8;
    assign CHOR05_n = CHOR05_n_U16004_10 & CHOR05_n_U16044_2 & CHOR05_n_U17003_10 & CHOR05_n_U17041_8 & CHOR05_n_U24011_10;
    assign CHOR06_n = CHOR06_n_U16004_12 & CHOR06_n_U16044_4 & CHOR06_n_U17003_12 & CHOR06_n_U17041_10 & CHOR06_n_U24011_12;
    assign CHOR07_n = CHOR07_n_U16021_2 & CHOR07_n_U16044_6 & CHOR07_n_U17012_2 & CHOR07_n_U17027_12 & CHOR07_n_U24017_2;
    assign CHOR08_n = CHOR08_n_U16021_4 & CHOR08_n_U17012_4 & CHOR08_n_U17041_12 & CHOR08_n_U24017_4;
    assign CHOR09_n = CHOR09_n_U17012_6 & CHOR09_n_U17052_2 & CHOR09_n_U24017_6 & CHOR09_n_U24017_8;
    assign CHOR10_n = CHOR10_n_U17012_8 & CHOR10_n_U17052_4 & CHOR10_n_U24017_10 & CHOR10_n_U24017_12;
    assign CHOR11_n = CHOR11_n_U17012_10 & CHOR11_n_U17052_6 & CHOR11_n_U24021_2 & CHOR11_n_U24021_4;
    assign CHOR12_n = CHOR12_n_U17012_12 & CHOR12_n_U17052_8 & CHOR12_n_U24021_6;
    assign CHOR13_n = CHOR13_n_U17019_2 & CHOR13_n_U17052_10 & CHOR13_n_U24021_8;
    assign CHOR14_n = CHOR14_n_U17019_4 & CHOR14_n_U17052_12 & CHOR14_n_U24021_10;
    assign CHOR16_n = CHOR16_n_U17019_6 & CHOR16_n_U17061_2 & CHOR16_n_U24021_12;
    assign CI_n = CI_n_U4061_12 & CI_n_U5018_2 & CI_n_U5044_10 & CI_n_U6047_2;
    assign CO06 = CO06_U8041_2 & CO06_U8050_2;
    assign CO10 = CO10_U9041_2 & CO10_U9050_2;
    assign CO14 = CO14_U10041_2 & CO14_U10050_2;
    assign G01_n = G01_n_U8013_6 & G01_n_U8013_8;
    assign G05_n = G05_n_U9013_6 & G05_n_U9013_8;
    assign G06_n = G06_n_U9028_10 & G06_n_U9028_12;
    assign G07_n = G07_n_U9050_6 & G07_n_U9050_8;
    assign G09_n = G09_n_U10013_6 & G09_n_U10013_8;
    assign G10_n = G10_n_U10028_10 & G10_n_U10028_12;
    assign G11_n = G11_n_U10050_6 & G11_n_U10050_8;
    assign G13_n = G13_n_U11013_6 & G13_n_U11013_8;
    assign G14_n = G14_n_U11028_10 & G14_n_U11028_12;
    assign G15_n = G15_n_U11050_6 & G15_n_U11050_8;
    assign GTONE = GTONE_U24029_2 & GTONE_U24029_4;
    assign INHPLS = INHPLS_U12016_10 & INHPLS_U12016_12;
    assign L01_n = L01_n_U8007_6;
    assign L02_n = L02_n_U8013_12;
    assign L04_n = L04_n_U8050_12;
    assign L08_n = L08_n_U9050_12;
    assign L12_n = L12_n_U10050_12;
    assign L15_n = L15_n_U11041_6;
    assign L16_n = L16_n_U4063_8 & L16_n_U11050_12;
    assign MONEX_n = MONEX_n_U5005_2 & MONEX_n_U6029_6;
    assign PALE = PALE_U12027_2 & PALE_U12027_4;
    assign R1C_n = R1C_n_U4063_10 & R1C_n_U6029_12;
    assign RA_n = RA_n_U4039_10 & RA_n_U4045_8 & RA_n_U5005_8 & RA_n_U5024_4 & RA_n_U5039_12;
    assign RB1_n = RB1_n_U4063_6 & RB1_n_U6029_10;
    assign RB_n = RB_n_U4039_2 & RB_n_U4061_10 & RB_n_U5005_6 & RB_n_U5018_10 & RB_n_U5049_2 & RB_n_U6004_8 & RB_n_U6037_8;
    assign RC_n = RC_n_U4039_4 & RC_n_U4061_8 & RC_n_U5012_8 & RC_n_U5024_10 & RC_n_U5049_10 & RC_n_U6047_6 & RC_n_U6052_8;
    assign RELPLS = RELPLS_U12016_6 & RELPLS_U12016_8;
    assign RG_n = RG_n_U5012_6 & RG_n_U5044_2 & RG_n_U5044_4 & RG_n_U5059_10 & RG_n_U6014_8;
    assign RL01_n = RL01_n_U8007_4 & RL01_n_U8007_10 & RL01_n_U8007_12 & RL01_n_U8013_4 & RL01_n_U15039_12;
    assign RL02_n = RL02_n_U8013_10 & RL02_n_U8028_2 & RL02_n_U8028_6 & RL02_n_U8028_8 & RL02_n_U15039_10;
    assign RL03_n = RL03_n_U8041_4 & RL03_n_U8041_10 & RL03_n_U8041_12 & RL03_n_U8050_4 & RL03_n_U15039_4;
    assign RL04_n = RL04_n_U8050_10 & RL04_n_U8061_2 & RL04_n_U8061_6 & RL04_n_U8061_8 & RL04_n_U15039_6;
    assign RL05_n = RL05_n_U9007_4 & RL05_n_U9007_10 & RL05_n_U9007_12 & RL05_n_U9013_4 & RL05_n_U15039_8;
    assign RL06_n = RL06_n_U9013_10 & RL06_n_U9028_2 & RL06_n_U9028_6 & RL06_n_U9028_8 & RL06_n_U15016_6;
    assign RL09_n = RL09_n_U10007_4 & RL09_n_U10007_10 & RL09_n_U10007_12 & RL09_n_U10013_4 & RL09_n_U15016_4;
    assign RL10_n = RL10_n_U10013_10 & RL10_n_U10028_2 & RL10_n_U10028_6 & RL10_n_U10028_8 & RL10_n_U15016_2;
    assign RL11_n = RL11_n_U10041_4 & RL11_n_U10041_10 & RL11_n_U10041_12 & RL11_n_U10050_4 & RL11_n_U15004_12;
    assign RL12_n = RL12_n_U10050_10 & RL12_n_U10061_2 & RL12_n_U10061_6 & RL12_n_U10061_8 & RL12_n_U15004_10;
    assign RL13_n = RL13_n_U11007_4 & RL13_n_U11007_10 & RL13_n_U11007_12 & RL13_n_U11013_4 & RL13_n_U15004_8;
    assign RL14_n = RL14_n_U11013_10 & RL14_n_U11028_2 & RL14_n_U11028_6 & RL14_n_U11028_8 & RL14_n_U15004_6;
    assign RL15_n = RL15_n_U11041_4 & RL15_n_U11041_10 & RL15_n_U11041_12 & RL15_n_U11050_4 & RL15_n_U15004_4;
    assign RL16_n = RL16_n_U11050_10 & RL16_n_U11061_2 & RL16_n_U11061_6 & RL16_n_U11061_8 & RL16_n_U15004_2;
    assign RL_n = RL_n_U5005_12 & RL_n_U5039_10;
    assign RPTSET = RPTSET_U3011_2 & RPTSET_U3011_4 & RPTSET_U3011_6 & RPTSET_U6052_4;
    assign RU_n = RU_n_U5024_2 & RU_n_U5059_4 & RU_n_U5059_6 & RU_n_U6014_12 & RU_n_U6037_2 & RU_n_U6052_6;
    assign RZ_n = RZ_n_U5005_4 & RZ_n_U5018_4 & RZ_n_U5049_4 & RZ_n_U6052_2;
    assign SCAD = SCAD_U5049_6 & SCAD_U5049_8;
    assign ST2_n = ST2_n_U5024_6 & ST2_n_U6047_12;
    assign TMZ_n = TMZ_n_U4045_12 & TMZ_n_U5012_2 & TMZ_n_U5065_6;
    assign TOV_n = TOV_n_U5059_2 & TOV_n_U6019_4;
    assign TSGN_n = TSGN_n_U4063_2 & TSGN_n_U4063_4 & TSGN_n_U5059_12 & TSGN_n_U5065_10;
    assign WA_n = WA_n_U5005_10 & WA_n_U5024_12 & WA_n_U5056_6 & WA_n_U6029_8 & WA_n_U6047_4;
    assign WB_n = WB_n_U5018_12 & WB_n_U5039_2 & WB_n_U5039_4 & WB_n_U5059_8 & WB_n_U6014_10;
    assign WG_n = WG_n_U4039_12 & WG_n_U4045_2 & WG_n_U4045_10 & WG_n_U5012_4 & WG_n_U6019_8 & WG_n_U6037_6;
    assign WL_n = WL_n_U4061_6 & WL_n_U5065_4 & WL_n_U6014_6;
    assign WSC_n = WSC_n_U6019_6 & WSC_n_U6037_4;
    assign WS_n = WS_n_U5034_12 & WS_n_U6041_8;
    assign WY12_n = WY12_n_U5018_6 & WY12_n_U5044_12;
    assign WYD_n = WYD_n_U5065_8 & WYD_n_U6004_10;
    assign WY_n = WY_n_U4061_2 & WY_n_U4061_4 & WY_n_U5012_12 & WY_n_U5024_8 & WY_n_U5044_6 & WY_n_U6004_12;
    assign WZ_n = WZ_n_U5018_8 & WZ_n_U5056_12 & WZ_n_U6019_2;
    assign Z15_n = Z15_n_U5065_2 & Z15_n_U11041_8;
    assign Z16_n = Z16_n_U5056_4 & Z16_n_U11061_4;
    assign __A02_1__Q2A = __A02_1__Q2A_U2148_4;
    assign __A02_3__T12SET = __A02_3__T12SET_U2038_2 & __A02_3__T12SET_U2038_4 & __A02_3__T12SET_U2038_6 & __A02_3__T12SET_U2038_8;
    assign __A02_NET_151 = __A02_NET_151_U2120_2 & __A02_NET_151_U2120_4;
    assign __A03_2__IC13_n = __A03_2__IC13_n_U3011_8 & __A03_2__IC13_n_U3011_10;
    assign __A04_1__SGUM = __A04_1__SGUM_U4003_10 & __A04_1__SGUM_U4003_12;
    assign __A04_NET_193 = __A04_NET_193_U4023_6 & __A04_NET_193_U4023_8;
    assign __A04_NET_204 = __A04_NET_204_U4023_10 & __A04_NET_204_U4023_12 & __A04_NET_204_U4029_2 & __A04_NET_204_U4029_4 & __A04_NET_204_U4029_6;
    assign __A04_NET_208 = __A04_NET_208_U4029_8 & __A04_NET_208_U4029_10;
    assign __A04_NET_215 = __A04_NET_215_U4023_2 & __A04_NET_215_U4023_4;
    assign __A04_NET_236 = __A04_NET_236_U4003_6 & __A04_NET_236_U4003_8;
    assign __A04_NET_249 = __A04_NET_249_U4003_2 & __A04_NET_249_U4003_4;
    assign __A04_NET_279 = __A04_NET_279_U4045_4 & __A04_NET_279_U4045_6;
    assign __A05_NET_260 = __A05_NET_260_U5049_12 & __A05_NET_260_U5056_2;
    assign __A05_NET_267 = __A05_NET_267_U5056_8 & __A05_NET_267_U5056_10;
    assign __A05_NET_282 = __A05_NET_282_U5034_8 & __A05_NET_282_U5034_10;
    assign __A05_NET_285 = __A05_NET_285_U5039_6 & __A05_NET_285_U5039_8;
    assign __A06_NET_186 = __A06_NET_186_U6041_10 & __A06_NET_186_U6041_12;
    assign __A06_NET_199 = __A06_NET_199_U6041_4 & __A06_NET_199_U6041_6;
    assign __A06_NET_203 = __A06_NET_203_U6019_10 & __A06_NET_203_U6019_12;
    assign __A06_NET_220 = __A06_NET_220_U6047_8 & __A06_NET_220_U6047_10;
    assign __A06_NET_241 = __A06_NET_241_U6029_2 & __A06_NET_241_U6029_4;
    assign __A06_NET_272 = __A06_NET_272_U6004_2 & __A06_NET_272_U6004_4;
    assign __A06_NET_320 = __A06_NET_320_U6014_2 & __A06_NET_320_U6014_4;
    assign __A07_NET_158 = __A07_NET_158_U7007_2 & __A07_NET_158_U7007_4;
    assign __A08_1___G2_n = __A08_1___G2_n_U8028_10 & __A08_1___G2_n_U8028_12;
    assign __A08_1___Z1_n = __A08_1___Z1_n_U8007_8;
    assign __A08_1___Z2_n = __A08_1___Z2_n_U8028_4;
    assign __A08_2___G1_n = __A08_2___G1_n_U8050_6 & __A08_2___G1_n_U8050_8;
    assign __A08_2___Z1_n = __A08_2___Z1_n_U8041_8;
    assign __A08_2___Z2_n = __A08_2___Z2_n_U8061_4;
    assign __A09_1___Z1_n = __A09_1___Z1_n_U9007_8;
    assign __A09_1___Z2_n = __A09_1___Z2_n_U9028_4;
    assign __A09_2___RL1_n = __A09_2___RL1_n_U9041_4 & __A09_2___RL1_n_U9041_10 & __A09_2___RL1_n_U9041_12 & __A09_2___RL1_n_U9050_4;
    assign __A09_2___RL2_n = __A09_2___RL2_n_U9050_10 & __A09_2___RL2_n_U9061_2 & __A09_2___RL2_n_U9061_6 & __A09_2___RL2_n_U9061_8;
    assign __A09_2___Z1_n = __A09_2___Z1_n_U9041_8;
    assign __A09_2___Z2_n = __A09_2___Z2_n_U9061_4;
    assign __A10_1___Z1_n = __A10_1___Z1_n_U10007_8;
    assign __A10_1___Z2_n = __A10_1___Z2_n_U10028_4;
    assign __A10_2___Z1_n = __A10_2___Z1_n_U10041_8;
    assign __A10_2___Z2_n = __A10_2___Z2_n_U10061_4;
    assign __A11_1___Z1_n = __A11_1___Z1_n_U11007_8;
    assign __A11_1___Z2_n = __A11_1___Z2_n_U11028_4;
    assign __A11_2___CO_OUT = __A11_2___CO_OUT_U11041_2 & __A11_2___CO_OUT_U11050_2;
    assign __A12_1__GNZRO = __A12_1__GNZRO_U12016_2 & __A12_1__GNZRO_U12016_4;
    assign __A13_1__CKTAL_n = __A13_1__CKTAL_n_U13006_2 & __A13_1__CKTAL_n_U13006_4;
    assign __A13_NET_179 = __A13_NET_179_U13121_2 & __A13_NET_179_U13121_4;
    assign __A13_NET_277 = __A13_NET_277_U13006_6 & __A13_NET_277_U13006_8 & __A13_NET_277_U13006_10 & __A13_NET_277_U13006_12 & __A13_NET_277_U13036_2 & __A13_NET_277_U13036_4 & __A13_NET_277_U13036_6 & __A13_NET_277_U13036_12 & __A13_NET_277_U13051_2 & __A13_NET_277_U13051_4 & __A13_NET_277_U13051_6;
    assign __A13_NET_307 = __A13_NET_307_U13036_8 & __A13_NET_307_U13036_10;
    assign __A14_1__ERAS = __A14_1__ERAS_U14014_10 & __A14_1__ERAS_U14014_12;
    assign __A14_1__SBFSET = __A14_1__SBFSET_U14014_2 & __A14_1__SBFSET_U14014_4;
    assign __A14_1__TPGE = __A14_1__TPGE_U14033_2 & __A14_1__TPGE_U14033_4;
    assign __A14_1__TPGF = __A14_1__TPGF_U14014_6 & __A14_1__TPGF_U14014_8;
    assign __A15_NET_229 = __A15_NET_229_U15016_8 & __A15_NET_229_U15016_10;
    assign __A15_NET_232 = __A15_NET_232_U15016_12 & __A15_NET_232_U15039_2;
    assign __A17_NET_176 = __A17_NET_176_U17019_8 & __A17_NET_176_U17019_10;
    assign __A17_NET_183 = __A17_NET_183_U17019_12 & __A17_NET_183_U17027_2;
    assign __A17_NET_220 = __A17_NET_220_U17027_4 & __A17_NET_220_U17027_6 & __A17_NET_220_U17027_8;
    assign __A18_2__CNTOF9 = __A18_2__CNTOF9_U18007_10 & __A18_2__CNTOF9_U18007_12;
    assign __A18_NET_116 = __A18_NET_116_U18007_2 & __A18_NET_116_U18007_4;
    assign __A18_NET_99 = __A18_NET_99_U18007_6 & __A18_NET_99_U18007_8;
    assign __A21_1__32004K = __A21_1__32004K_U21010_2 & __A21_1__32004K_U21010_4;
    assign __A21_NET_141 = __A21_NET_141_U21023_2 & __A21_NET_141_U21023_4 & __A21_NET_141_U21023_6;
    assign __A21_NET_145 = __A21_NET_145_U21023_8 & __A21_NET_145_U21023_10;
    assign __A21_NET_146 = __A21_NET_146_U21010_10 & __A21_NET_146_U21010_12;
    assign __A21_NET_147 = __A21_NET_147_U21006_6 & __A21_NET_147_U21006_8 & __A21_NET_147_U21006_10 & __A21_NET_147_U21006_12;
    assign __A21_NET_152 = __A21_NET_152_U21002_2 & __A21_NET_152_U21002_4 & __A21_NET_152_U21002_6 & __A21_NET_152_U21002_8;
    assign __A21_NET_153 = __A21_NET_153_U21002_10 & __A21_NET_153_U21002_12 & __A21_NET_153_U21006_2 & __A21_NET_153_U21006_4;
    assign __A21_NET_159 = __A21_NET_159_U21023_12 & __A21_NET_159_U21027_2;
    assign __A21_NET_162 = __A21_NET_162_U21027_4 & __A21_NET_162_U21027_6;
    assign __A21_NET_173 = __A21_NET_173_U21010_6 & __A21_NET_173_U21010_8;
    assign __A21_NET_187 = __A21_NET_187_U21014_2 & __A21_NET_187_U21014_4 & __A21_NET_187_U21014_6;
    assign __A21_NET_229 = __A21_NET_229_U21014_8 & __A21_NET_229_U21014_10 & __A21_NET_229_U21014_12;
    assign __A22_1__DATA_n = __A22_1__DATA_n_U22028_2 & __A22_1__DATA_n_U22028_4 & __A22_1__DATA_n_U22028_6 & __A22_1__DATA_n_U22028_8 & __A22_1__DATA_n_U22028_10 & __A22_1__DATA_n_U22028_12 & __A22_1__DATA_n_U22057_2 & __A22_1__DATA_n_U22057_4 & __A22_1__DATA_n_U22057_6;
    assign __A23_NET_174 = __A23_NET_174_U23002_6 & __A23_NET_174_U23002_8;
    assign __A23_NET_185 = __A23_NET_185_U23002_2 & __A23_NET_185_U23002_4;
    assign __CO04 = __CO04_U8007_2 & __CO04_U8013_2;
    assign __CO08 = __CO08_U9007_2 & __CO08_U9013_2;
    assign __CO12 = __CO12_U10007_2 & __CO12_U10013_2;
    assign __CO16 = __CO16_U11007_2 & __CO16_U11013_2;
    assign __G04_n = __G04_n_U8061_10 & __G04_n_U8061_12;
    assign __G08_n = __G08_n_U9061_10 & __G08_n_U9061_12;
    assign __G12_n = __G12_n_U10061_10 & __G12_n_U10061_12;
    assign __G16_n = __G16_n_U11061_10 & __G16_n_U11061_12;
    assign __L03_n = __L03_n_U8041_6;
    assign __L05_n = __L05_n_U9007_6;
    assign __L06_n = __L06_n_U9013_12;
    assign __L07_n = __L07_n_U9041_6;
    assign __L09_n = __L09_n_U10007_6;
    assign __L10_n = __L10_n_U10013_12;
    assign __L11_n = __L11_n_U10041_6;
    assign __L13_n = __L13_n_U11007_6;
    assign __L14_n = __L14_n_U11013_12;
    assign n5XP11 = n5XP11_U4039_6 & n5XP11_U4039_8;
    assign n8PP4 = n8PP4_U4063_12 & n8PP4_U6037_10 & n8PP4_U6037_12 & n8PP4_U6041_2;
    assign SA01 = GND | SA01_U31001_29 | SA01_U31023_16 | SA01_U31025_7;
    assign SA02 = GND | SA02_U31001_31 | SA02_U31023_14 | SA02_U31025_8;
    assign SA03 = GND | SA03_U31001_33 | SA03_U31023_12 | SA03_U31025_9;
    assign SA04 = GND | SA04_U31001_35 | SA04_U31023_9 | SA04_U31025_10;
    assign SA05 = GND | SA05_U31001_38 | SA05_U31023_7 | SA05_U31025_13;
    assign SA06 = GND | SA06_U31001_40 | SA06_U31023_5 | SA06_U31025_14;
    assign SA07 = GND | SA07_U31001_42 | SA07_U31023_3 | SA07_U31025_15;
    assign SA08 = GND | SA08_U31001_44 | SA08_U31024_18 | SA08_U31025_16;
    assign SA09 = GND | SA09_U31001_30 | SA09_U31024_16 | SA09_U31025_29;
    assign SA10 = GND | SA10_U31001_32 | SA10_U31024_14 | SA10_U31025_30;
    assign SA11 = GND | SA11_U31001_34 | SA11_U31024_12 | SA11_U31025_31;
    assign SA12 = GND | SA12_U31001_36 | SA12_U31024_9 | SA12_U31025_32;
    assign SA13 = GND | SA13_U31001_39 | SA13_U31024_7 | SA13_U31025_35;
    assign SA14 = GND | SA14_U31001_41 | SA14_U31024_5 | SA14_U31025_36;
    assign SA16 = GND | SA16_U31001_45 | SA16_U31024_3 | SA16_U31025_38;
    assign SAP = GND | SAP_U31001_43 | SAP_U31023_18 | SAP_U31025_37;
endmodule
`default_nettype wire
